module ripple_carry_adder_routing (cin,
    clk,
    cout,
    overflow,
    a,
    b,
    sum);
 input cin;
 input clk;
 output cout;
 output overflow;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire \bit_adder[0].FA.sum ;
 wire \bit_adder[10].FA.sum ;
 wire \bit_adder[11].FA.sum ;
 wire \bit_adder[12].FA.sum ;
 wire \bit_adder[13].FA.sum ;
 wire \bit_adder[14].FA.sum ;
 wire \bit_adder[15].FA.sum ;
 wire \bit_adder[16].FA.sum ;
 wire \bit_adder[17].FA.sum ;
 wire \bit_adder[18].FA.sum ;
 wire \bit_adder[19].FA.sum ;
 wire \bit_adder[1].FA.sum ;
 wire \bit_adder[20].FA.sum ;
 wire \bit_adder[21].FA.sum ;
 wire \bit_adder[22].FA.sum ;
 wire \bit_adder[23].FA.sum ;
 wire \bit_adder[24].FA.sum ;
 wire \bit_adder[25].FA.sum ;
 wire \bit_adder[26].FA.sum ;
 wire \bit_adder[27].FA.sum ;
 wire \bit_adder[28].FA.sum ;
 wire \bit_adder[29].FA.sum ;
 wire \bit_adder[2].FA.sum ;
 wire \bit_adder[30].FA.sum ;
 wire \bit_adder[31].FA.sum ;
 wire \bit_adder[3].FA.sum ;
 wire \bit_adder[4].FA.sum ;
 wire \bit_adder[5].FA.sum ;
 wire \bit_adder[6].FA.sum ;
 wire \bit_adder[7].FA.sum ;
 wire \bit_adder[8].FA.sum ;
 wire \bit_adder[9].FA.sum ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__inv_2 _216_ (.A(net56),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _217_ (.A(net24),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _218_ (.A(net53),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _219_ (.A(net21),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _220_ (.A(net51),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _221_ (.A(net19),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _222_ (.A(net48),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _223_ (.A(net16),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _224_ (.A(net46),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _225_ (.A(net14),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _226_ (.A(net45),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _227_ (.A(net13),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _228_ (.A(net42),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _229_ (.A(net10),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _230_ (.A(net40),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _231_ (.A(net8),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _232_ (.A(net39),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _233_ (.A(net7),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _234_ (.A(net37),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _235_ (.A(net5),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _236_ (.A(net35),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _237_ (.A(net3),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _238_ (.A(net34),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(net2),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(net63),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _241_ (.A(net31),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _242_ (.A(net61),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _243_ (.A(net29),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _244_ (.A(net59),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _245_ (.A(net27),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _246_ (.A(net55),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _247_ (.A(net23),
    .Y(_031_));
 sky130_fd_sc_hd__nor2_1 _248_ (.A(net57),
    .B(net25),
    .Y(_032_));
 sky130_fd_sc_hd__or2_1 _249_ (.A(net57),
    .B(net25),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _250_ (.A(net57),
    .B(net25),
    .X(_034_));
 sky130_fd_sc_hd__nand2_1 _251_ (.A(net57),
    .B(net25),
    .Y(_035_));
 sky130_fd_sc_hd__or2_1 _252_ (.A(net56),
    .B(net24),
    .X(_036_));
 sky130_fd_sc_hd__nor2_1 _253_ (.A(_000_),
    .B(_001_),
    .Y(_037_));
 sky130_fd_sc_hd__nand2_1 _254_ (.A(net56),
    .B(net24),
    .Y(_038_));
 sky130_fd_sc_hd__or2_1 _255_ (.A(net54),
    .B(net22),
    .X(_039_));
 sky130_fd_sc_hd__nand2_2 _256_ (.A(net54),
    .B(net22),
    .Y(_040_));
 sky130_fd_sc_hd__or2_1 _257_ (.A(net53),
    .B(net21),
    .X(_041_));
 sky130_fd_sc_hd__nand2_1 _258_ (.A(net53),
    .B(net21),
    .Y(_042_));
 sky130_fd_sc_hd__or2_1 _259_ (.A(net52),
    .B(net20),
    .X(_043_));
 sky130_fd_sc_hd__nand2_2 _260_ (.A(net52),
    .B(net20),
    .Y(_044_));
 sky130_fd_sc_hd__or2_1 _261_ (.A(net51),
    .B(net19),
    .X(_045_));
 sky130_fd_sc_hd__nand2_1 _262_ (.A(net51),
    .B(net19),
    .Y(_046_));
 sky130_fd_sc_hd__or2_1 _263_ (.A(net50),
    .B(net18),
    .X(_047_));
 sky130_fd_sc_hd__nand2_1 _264_ (.A(net50),
    .B(net18),
    .Y(_048_));
 sky130_fd_sc_hd__or2_1 _265_ (.A(net49),
    .B(net17),
    .X(_049_));
 sky130_fd_sc_hd__nand2_1 _266_ (.A(net49),
    .B(net17),
    .Y(_050_));
 sky130_fd_sc_hd__nand2_1 _267_ (.A(net48),
    .B(net16),
    .Y(_051_));
 sky130_fd_sc_hd__or2_1 _268_ (.A(net47),
    .B(net15),
    .X(_052_));
 sky130_fd_sc_hd__nand2_1 _269_ (.A(net47),
    .B(net15),
    .Y(_053_));
 sky130_fd_sc_hd__or2_1 _270_ (.A(net46),
    .B(net14),
    .X(_054_));
 sky130_fd_sc_hd__nand2_1 _271_ (.A(net46),
    .B(net14),
    .Y(_055_));
 sky130_fd_sc_hd__or2_1 _272_ (.A(net43),
    .B(net11),
    .X(_056_));
 sky130_fd_sc_hd__nand2_1 _273_ (.A(net43),
    .B(net11),
    .Y(_057_));
 sky130_fd_sc_hd__nor2_1 _274_ (.A(net42),
    .B(net10),
    .Y(_058_));
 sky130_fd_sc_hd__or2_1 _275_ (.A(net41),
    .B(net9),
    .X(_059_));
 sky130_fd_sc_hd__nand2_2 _276_ (.A(net41),
    .B(net9),
    .Y(_060_));
 sky130_fd_sc_hd__or2_1 _277_ (.A(net40),
    .B(net8),
    .X(_061_));
 sky130_fd_sc_hd__nand2_1 _278_ (.A(net40),
    .B(net8),
    .Y(_062_));
 sky130_fd_sc_hd__or2_2 _279_ (.A(net38),
    .B(net6),
    .X(_063_));
 sky130_fd_sc_hd__nand2_2 _280_ (.A(net38),
    .B(net6),
    .Y(_064_));
 sky130_fd_sc_hd__or2_1 _281_ (.A(net37),
    .B(net5),
    .X(_065_));
 sky130_fd_sc_hd__nor2_1 _282_ (.A(_018_),
    .B(_019_),
    .Y(_066_));
 sky130_fd_sc_hd__nand2_1 _283_ (.A(net37),
    .B(net5),
    .Y(_067_));
 sky130_fd_sc_hd__or2_1 _284_ (.A(net36),
    .B(net4),
    .X(_068_));
 sky130_fd_sc_hd__nand2_2 _285_ (.A(net36),
    .B(net4),
    .Y(_069_));
 sky130_fd_sc_hd__or2_1 _286_ (.A(net35),
    .B(net3),
    .X(_070_));
 sky130_fd_sc_hd__nand2_1 _287_ (.A(net35),
    .B(net3),
    .Y(_071_));
 sky130_fd_sc_hd__or2_1 _288_ (.A(net64),
    .B(net32),
    .X(_072_));
 sky130_fd_sc_hd__nand2_1 _289_ (.A(net64),
    .B(net32),
    .Y(_073_));
 sky130_fd_sc_hd__or2_1 _290_ (.A(net63),
    .B(net31),
    .X(_074_));
 sky130_fd_sc_hd__nand2_1 _291_ (.A(net63),
    .B(net31),
    .Y(_075_));
 sky130_fd_sc_hd__or2_1 _292_ (.A(net62),
    .B(net30),
    .X(_076_));
 sky130_fd_sc_hd__nand2_2 _293_ (.A(net62),
    .B(net30),
    .Y(_077_));
 sky130_fd_sc_hd__nand2_2 _294_ (.A(net60),
    .B(net28),
    .Y(_078_));
 sky130_fd_sc_hd__or2_1 _295_ (.A(net59),
    .B(net27),
    .X(_079_));
 sky130_fd_sc_hd__nor2_1 _296_ (.A(net58),
    .B(net26),
    .Y(_080_));
 sky130_fd_sc_hd__nand2_2 _297_ (.A(net58),
    .B(net26),
    .Y(_081_));
 sky130_fd_sc_hd__nand2_1 _298_ (.A(net44),
    .B(net12),
    .Y(_082_));
 sky130_fd_sc_hd__or2_1 _299_ (.A(net44),
    .B(net12),
    .X(_083_));
 sky130_fd_sc_hd__nand2_1 _300_ (.A(net1),
    .B(net65),
    .Y(_084_));
 sky130_fd_sc_hd__or2_1 _301_ (.A(net1),
    .B(net65),
    .X(_085_));
 sky130_fd_sc_hd__o21ai_1 _302_ (.A1(net1),
    .A2(net65),
    .B1(net33),
    .Y(_086_));
 sky130_fd_sc_hd__and2_1 _303_ (.A(_084_),
    .B(_086_),
    .X(_087_));
 sky130_fd_sc_hd__nand3_2 _304_ (.A(_082_),
    .B(_084_),
    .C(_086_),
    .Y(_088_));
 sky130_fd_sc_hd__o21ai_1 _305_ (.A1(net44),
    .A2(net12),
    .B1(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__o22a_1 _306_ (.A1(net55),
    .A2(net23),
    .B1(net44),
    .B2(net12),
    .X(_090_));
 sky130_fd_sc_hd__nand2_1 _307_ (.A(_088_),
    .B(_090_),
    .Y(_091_));
 sky130_fd_sc_hd__a22oi_4 _308_ (.A1(net55),
    .A2(net23),
    .B1(_088_),
    .B2(_090_),
    .Y(_092_));
 sky130_fd_sc_hd__o211ai_2 _309_ (.A1(_030_),
    .A2(_031_),
    .B1(_081_),
    .C1(_091_),
    .Y(_093_));
 sky130_fd_sc_hd__o21ai_1 _310_ (.A1(_080_),
    .A2(_092_),
    .B1(_081_),
    .Y(_094_));
 sky130_fd_sc_hd__o221ai_4 _311_ (.A1(_028_),
    .A2(_029_),
    .B1(_080_),
    .B2(_092_),
    .C1(_081_),
    .Y(_095_));
 sky130_fd_sc_hd__o221ai_4 _312_ (.A1(net59),
    .A2(net27),
    .B1(net58),
    .B2(net26),
    .C1(_093_),
    .Y(_096_));
 sky130_fd_sc_hd__o21ai_1 _313_ (.A1(net59),
    .A2(net27),
    .B1(_095_),
    .Y(_097_));
 sky130_fd_sc_hd__o211ai_4 _314_ (.A1(_028_),
    .A2(_029_),
    .B1(_078_),
    .C1(_096_),
    .Y(_098_));
 sky130_fd_sc_hd__o211ai_1 _315_ (.A1(net60),
    .A2(net28),
    .B1(_079_),
    .C1(_095_),
    .Y(_099_));
 sky130_fd_sc_hd__o21ai_1 _316_ (.A1(net60),
    .A2(net28),
    .B1(_098_),
    .Y(_100_));
 sky130_fd_sc_hd__o211ai_1 _317_ (.A1(_026_),
    .A2(_027_),
    .B1(_078_),
    .C1(_099_),
    .Y(_101_));
 sky130_fd_sc_hd__o221ai_4 _318_ (.A1(net61),
    .A2(net29),
    .B1(net60),
    .B2(net28),
    .C1(_098_),
    .Y(_102_));
 sky130_fd_sc_hd__o21ai_1 _319_ (.A1(net61),
    .A2(net29),
    .B1(_101_),
    .Y(_103_));
 sky130_fd_sc_hd__o211ai_4 _320_ (.A1(_026_),
    .A2(_027_),
    .B1(_077_),
    .C1(_102_),
    .Y(_104_));
 sky130_fd_sc_hd__o211ai_1 _321_ (.A1(net61),
    .A2(net29),
    .B1(_076_),
    .C1(_101_),
    .Y(_105_));
 sky130_fd_sc_hd__o21ai_1 _322_ (.A1(net62),
    .A2(net30),
    .B1(_104_),
    .Y(_106_));
 sky130_fd_sc_hd__o211ai_1 _323_ (.A1(_024_),
    .A2(_025_),
    .B1(_077_),
    .C1(_105_),
    .Y(_107_));
 sky130_fd_sc_hd__o221ai_4 _324_ (.A1(net63),
    .A2(net31),
    .B1(net62),
    .B2(net30),
    .C1(_104_),
    .Y(_108_));
 sky130_fd_sc_hd__o21ai_1 _325_ (.A1(_024_),
    .A2(_025_),
    .B1(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__o211ai_2 _326_ (.A1(_024_),
    .A2(_025_),
    .B1(_073_),
    .C1(_108_),
    .Y(_110_));
 sky130_fd_sc_hd__o211ai_1 _327_ (.A1(net63),
    .A2(net31),
    .B1(_072_),
    .C1(_107_),
    .Y(_111_));
 sky130_fd_sc_hd__o21ai_1 _328_ (.A1(net64),
    .A2(net32),
    .B1(_110_),
    .Y(_112_));
 sky130_fd_sc_hd__o211ai_2 _329_ (.A1(_022_),
    .A2(_023_),
    .B1(_073_),
    .C1(_111_),
    .Y(_113_));
 sky130_fd_sc_hd__o221ai_2 _330_ (.A1(net34),
    .A2(net2),
    .B1(net64),
    .B2(net32),
    .C1(_110_),
    .Y(_114_));
 sky130_fd_sc_hd__o21ai_1 _331_ (.A1(net34),
    .A2(net2),
    .B1(_113_),
    .Y(_115_));
 sky130_fd_sc_hd__o221ai_2 _332_ (.A1(_020_),
    .A2(_021_),
    .B1(_022_),
    .B2(_023_),
    .C1(_114_),
    .Y(_116_));
 sky130_fd_sc_hd__o211ai_4 _333_ (.A1(net34),
    .A2(net2),
    .B1(_070_),
    .C1(_113_),
    .Y(_117_));
 sky130_fd_sc_hd__o21ai_1 _334_ (.A1(_020_),
    .A2(_021_),
    .B1(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__o211ai_4 _335_ (.A1(_020_),
    .A2(_021_),
    .B1(_069_),
    .C1(_117_),
    .Y(_119_));
 sky130_fd_sc_hd__o221ai_2 _336_ (.A1(net36),
    .A2(net4),
    .B1(net35),
    .B2(net3),
    .C1(_116_),
    .Y(_120_));
 sky130_fd_sc_hd__o21ai_1 _337_ (.A1(net36),
    .A2(net4),
    .B1(_119_),
    .Y(_121_));
 sky130_fd_sc_hd__o211ai_2 _338_ (.A1(_018_),
    .A2(_019_),
    .B1(_069_),
    .C1(_120_),
    .Y(_122_));
 sky130_fd_sc_hd__o221a_1 _339_ (.A1(net37),
    .A2(net5),
    .B1(net36),
    .B2(net4),
    .C1(_119_),
    .X(_123_));
 sky130_fd_sc_hd__o211ai_2 _340_ (.A1(net36),
    .A2(net4),
    .B1(_065_),
    .C1(_119_),
    .Y(_124_));
 sky130_fd_sc_hd__o211ai_4 _341_ (.A1(_018_),
    .A2(_019_),
    .B1(_064_),
    .C1(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__o221ai_4 _342_ (.A1(net38),
    .A2(net6),
    .B1(net37),
    .B2(net5),
    .C1(_122_),
    .Y(_126_));
 sky130_fd_sc_hd__o21ai_4 _343_ (.A1(net38),
    .A2(net6),
    .B1(_125_),
    .Y(_127_));
 sky130_fd_sc_hd__o211ai_2 _344_ (.A1(_016_),
    .A2(_017_),
    .B1(_064_),
    .C1(_126_),
    .Y(_128_));
 sky130_fd_sc_hd__o211ai_4 _345_ (.A1(net39),
    .A2(net7),
    .B1(_063_),
    .C1(_125_),
    .Y(_129_));
 sky130_fd_sc_hd__o21ai_4 _346_ (.A1(_016_),
    .A2(_017_),
    .B1(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__o211ai_4 _347_ (.A1(_016_),
    .A2(_017_),
    .B1(_062_),
    .C1(_129_),
    .Y(_131_));
 sky130_fd_sc_hd__o221ai_4 _348_ (.A1(net40),
    .A2(net8),
    .B1(net39),
    .B2(net7),
    .C1(_128_),
    .Y(_132_));
 sky130_fd_sc_hd__o21ai_1 _349_ (.A1(_014_),
    .A2(_015_),
    .B1(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__o211ai_4 _350_ (.A1(_014_),
    .A2(_015_),
    .B1(_060_),
    .C1(_132_),
    .Y(_134_));
 sky130_fd_sc_hd__o211ai_2 _351_ (.A1(net40),
    .A2(net8),
    .B1(_059_),
    .C1(_131_),
    .Y(_135_));
 sky130_fd_sc_hd__o21ai_1 _352_ (.A1(net41),
    .A2(net9),
    .B1(_134_),
    .Y(_136_));
 sky130_fd_sc_hd__o211ai_1 _353_ (.A1(_012_),
    .A2(_013_),
    .B1(_060_),
    .C1(_135_),
    .Y(_137_));
 sky130_fd_sc_hd__o221ai_4 _354_ (.A1(net42),
    .A2(net10),
    .B1(net41),
    .B2(net9),
    .C1(_134_),
    .Y(_138_));
 sky130_fd_sc_hd__o21ai_1 _355_ (.A1(_012_),
    .A2(_013_),
    .B1(_138_),
    .Y(_139_));
 sky130_fd_sc_hd__o21ai_1 _356_ (.A1(net42),
    .A2(net10),
    .B1(_137_),
    .Y(_140_));
 sky130_fd_sc_hd__o211ai_4 _357_ (.A1(_012_),
    .A2(_013_),
    .B1(_057_),
    .C1(_138_),
    .Y(_141_));
 sky130_fd_sc_hd__o211ai_1 _358_ (.A1(net42),
    .A2(net10),
    .B1(_056_),
    .C1(_137_),
    .Y(_142_));
 sky130_fd_sc_hd__o21ai_1 _359_ (.A1(net43),
    .A2(net11),
    .B1(_141_),
    .Y(_143_));
 sky130_fd_sc_hd__o211ai_1 _360_ (.A1(_010_),
    .A2(_011_),
    .B1(_057_),
    .C1(_142_),
    .Y(_144_));
 sky130_fd_sc_hd__o221ai_4 _361_ (.A1(net45),
    .A2(net13),
    .B1(net43),
    .B2(net11),
    .C1(_141_),
    .Y(_145_));
 sky130_fd_sc_hd__o21ai_1 _362_ (.A1(_010_),
    .A2(_011_),
    .B1(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__o221ai_2 _363_ (.A1(_008_),
    .A2(_009_),
    .B1(_010_),
    .B2(_011_),
    .C1(_145_),
    .Y(_147_));
 sky130_fd_sc_hd__o211ai_1 _364_ (.A1(net45),
    .A2(net13),
    .B1(_054_),
    .C1(_144_),
    .Y(_148_));
 sky130_fd_sc_hd__o21ai_1 _365_ (.A1(_008_),
    .A2(_009_),
    .B1(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__o211ai_1 _366_ (.A1(_008_),
    .A2(_009_),
    .B1(_053_),
    .C1(_148_),
    .Y(_150_));
 sky130_fd_sc_hd__o221ai_2 _367_ (.A1(net47),
    .A2(net15),
    .B1(net46),
    .B2(net14),
    .C1(_147_),
    .Y(_151_));
 sky130_fd_sc_hd__o21ai_1 _368_ (.A1(net47),
    .A2(net15),
    .B1(_150_),
    .Y(_152_));
 sky130_fd_sc_hd__o211ai_2 _369_ (.A1(_006_),
    .A2(_007_),
    .B1(_053_),
    .C1(_151_),
    .Y(_153_));
 sky130_fd_sc_hd__o211ai_1 _370_ (.A1(net48),
    .A2(net16),
    .B1(_052_),
    .C1(_150_),
    .Y(_154_));
 sky130_fd_sc_hd__o21ai_1 _371_ (.A1(net48),
    .A2(net16),
    .B1(_153_),
    .Y(_155_));
 sky130_fd_sc_hd__o211ai_1 _372_ (.A1(_006_),
    .A2(_007_),
    .B1(_050_),
    .C1(_154_),
    .Y(_156_));
 sky130_fd_sc_hd__o221ai_2 _373_ (.A1(net49),
    .A2(net17),
    .B1(net48),
    .B2(net16),
    .C1(_153_),
    .Y(_157_));
 sky130_fd_sc_hd__o21ai_1 _374_ (.A1(net49),
    .A2(net17),
    .B1(_156_),
    .Y(_158_));
 sky130_fd_sc_hd__nand3_2 _375_ (.A(_048_),
    .B(_050_),
    .C(_157_),
    .Y(_159_));
 sky130_fd_sc_hd__o211ai_1 _376_ (.A1(net49),
    .A2(net17),
    .B1(_047_),
    .C1(_156_),
    .Y(_160_));
 sky130_fd_sc_hd__o211ai_1 _377_ (.A1(_004_),
    .A2(_005_),
    .B1(_048_),
    .C1(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__o221ai_4 _378_ (.A1(net51),
    .A2(net19),
    .B1(net50),
    .B2(net18),
    .C1(_159_),
    .Y(_162_));
 sky130_fd_sc_hd__o21ai_1 _379_ (.A1(_004_),
    .A2(_005_),
    .B1(_162_),
    .Y(_163_));
 sky130_fd_sc_hd__o211ai_2 _380_ (.A1(_004_),
    .A2(_005_),
    .B1(_044_),
    .C1(_162_),
    .Y(_164_));
 sky130_fd_sc_hd__o211ai_2 _381_ (.A1(net51),
    .A2(net19),
    .B1(_043_),
    .C1(_161_),
    .Y(_165_));
 sky130_fd_sc_hd__o21ai_1 _382_ (.A1(net52),
    .A2(net20),
    .B1(_164_),
    .Y(_166_));
 sky130_fd_sc_hd__o211ai_4 _383_ (.A1(_002_),
    .A2(_003_),
    .B1(_044_),
    .C1(_165_),
    .Y(_167_));
 sky130_fd_sc_hd__o221ai_2 _384_ (.A1(net53),
    .A2(net21),
    .B1(net52),
    .B2(net20),
    .C1(_164_),
    .Y(_168_));
 sky130_fd_sc_hd__o211ai_2 _385_ (.A1(_002_),
    .A2(_003_),
    .B1(_040_),
    .C1(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__o211ai_4 _386_ (.A1(net53),
    .A2(net21),
    .B1(_039_),
    .C1(_167_),
    .Y(_170_));
 sky130_fd_sc_hd__o211ai_2 _387_ (.A1(_000_),
    .A2(_001_),
    .B1(_040_),
    .C1(_170_),
    .Y(_171_));
 sky130_fd_sc_hd__a2bb2oi_1 _388_ (.A1_N(net56),
    .A2_N(net24),
    .B1(_040_),
    .B2(_170_),
    .Y(_172_));
 sky130_fd_sc_hd__o221ai_2 _389_ (.A1(net56),
    .A2(net24),
    .B1(net54),
    .B2(net22),
    .C1(_169_),
    .Y(_173_));
 sky130_fd_sc_hd__o221ai_2 _390_ (.A1(net57),
    .A2(net25),
    .B1(net56),
    .B2(net24),
    .C1(_171_),
    .Y(_174_));
 sky130_fd_sc_hd__a31o_1 _391_ (.A1(_033_),
    .A2(_036_),
    .A3(_171_),
    .B1(_034_),
    .X(net66));
 sky130_fd_sc_hd__o31a_1 _392_ (.A1(_034_),
    .A2(_037_),
    .A3(_172_),
    .B1(_174_),
    .X(net67));
 sky130_fd_sc_hd__and3_1 _393_ (.A(net33),
    .B(net1),
    .C(net65),
    .X(_175_));
 sky130_fd_sc_hd__o22a_1 _394_ (.A1(_085_),
    .A2(net33),
    .B1(_175_),
    .B2(_087_),
    .X(\bit_adder[0].FA.sum ));
 sky130_fd_sc_hd__and3_1 _395_ (.A(_087_),
    .B(_083_),
    .C(_082_),
    .X(_176_));
 sky130_fd_sc_hd__a21oi_1 _396_ (.A1(_082_),
    .A2(_083_),
    .B1(_087_),
    .Y(_177_));
 sky130_fd_sc_hd__or2_1 _397_ (.A(_176_),
    .B(_177_),
    .X(\bit_adder[1].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _398_ (.A(net55),
    .B(net23),
    .X(_178_));
 sky130_fd_sc_hd__xnor2_1 _399_ (.A(_089_),
    .B(_178_),
    .Y(\bit_adder[2].FA.sum ));
 sky130_fd_sc_hd__and2b_1 _400_ (.A_N(_080_),
    .B(_081_),
    .X(_179_));
 sky130_fd_sc_hd__xnor2_1 _401_ (.A(_092_),
    .B(_179_),
    .Y(\bit_adder[3].FA.sum ));
 sky130_fd_sc_hd__and3_1 _402_ (.A(net59),
    .B(net27),
    .C(_094_),
    .X(_180_));
 sky130_fd_sc_hd__o22a_1 _403_ (.A1(_079_),
    .A2(_094_),
    .B1(_097_),
    .B2(_180_),
    .X(\bit_adder[4].FA.sum ));
 sky130_fd_sc_hd__a211o_1 _404_ (.A1(_079_),
    .A2(_095_),
    .B1(net60),
    .C1(net28),
    .X(_181_));
 sky130_fd_sc_hd__a2bb2o_1 _405_ (.A1_N(_078_),
    .A2_N(_097_),
    .B1(_100_),
    .B2(_181_),
    .X(\bit_adder[5].FA.sum ));
 sky130_fd_sc_hd__xnor2_1 _406_ (.A(net61),
    .B(net29),
    .Y(_182_));
 sky130_fd_sc_hd__xor2_1 _407_ (.A(_100_),
    .B(_182_),
    .X(\bit_adder[6].FA.sum ));
 sky130_fd_sc_hd__a21oi_1 _408_ (.A1(_076_),
    .A2(_077_),
    .B1(_103_),
    .Y(_183_));
 sky130_fd_sc_hd__and3_1 _409_ (.A(_076_),
    .B(_077_),
    .C(_103_),
    .X(_184_));
 sky130_fd_sc_hd__or2_1 _410_ (.A(_183_),
    .B(_184_),
    .X(\bit_adder[7].FA.sum ));
 sky130_fd_sc_hd__a21oi_1 _411_ (.A1(_074_),
    .A2(_075_),
    .B1(_106_),
    .Y(_185_));
 sky130_fd_sc_hd__and3_1 _412_ (.A(_074_),
    .B(_075_),
    .C(_106_),
    .X(_186_));
 sky130_fd_sc_hd__or2_1 _413_ (.A(_185_),
    .B(_186_),
    .X(\bit_adder[8].FA.sum ));
 sky130_fd_sc_hd__and3_1 _414_ (.A(net64),
    .B(net32),
    .C(_109_),
    .X(_187_));
 sky130_fd_sc_hd__o22a_1 _415_ (.A1(_072_),
    .A2(_109_),
    .B1(_112_),
    .B2(_187_),
    .X(\bit_adder[9].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _416_ (.A(net34),
    .B(net2),
    .X(_188_));
 sky130_fd_sc_hd__xnor2_1 _417_ (.A(_112_),
    .B(_188_),
    .Y(\bit_adder[10].FA.sum ));
 sky130_fd_sc_hd__nand2_1 _418_ (.A(_070_),
    .B(_071_),
    .Y(_189_));
 sky130_fd_sc_hd__xor2_1 _419_ (.A(_115_),
    .B(_189_),
    .X(\bit_adder[11].FA.sum ));
 sky130_fd_sc_hd__nand2_1 _420_ (.A(_068_),
    .B(_069_),
    .Y(_190_));
 sky130_fd_sc_hd__xnor2_1 _421_ (.A(_118_),
    .B(_190_),
    .Y(\bit_adder[12].FA.sum ));
 sky130_fd_sc_hd__nand2_1 _422_ (.A(_065_),
    .B(_067_),
    .Y(_191_));
 sky130_fd_sc_hd__xor2_1 _423_ (.A(_121_),
    .B(_191_),
    .X(\bit_adder[13].FA.sum ));
 sky130_fd_sc_hd__and4_1 _424_ (.A(_122_),
    .B(net6),
    .C(net38),
    .D(_065_),
    .X(_192_));
 sky130_fd_sc_hd__o32a_1 _425_ (.A1(_063_),
    .A2(_066_),
    .A3(_123_),
    .B1(_192_),
    .B2(_127_),
    .X(\bit_adder[14].FA.sum ));
 sky130_fd_sc_hd__xnor2_2 _426_ (.A(net39),
    .B(net7),
    .Y(_193_));
 sky130_fd_sc_hd__xor2_4 _427_ (.A(_127_),
    .B(_193_),
    .X(\bit_adder[15].FA.sum ));
 sky130_fd_sc_hd__nand2_2 _428_ (.A(_061_),
    .B(_062_),
    .Y(_194_));
 sky130_fd_sc_hd__xnor2_4 _429_ (.A(_130_),
    .B(_194_),
    .Y(\bit_adder[16].FA.sum ));
 sky130_fd_sc_hd__nand2_1 _430_ (.A(_059_),
    .B(_060_),
    .Y(_195_));
 sky130_fd_sc_hd__xnor2_1 _431_ (.A(_133_),
    .B(_195_),
    .Y(\bit_adder[17].FA.sum ));
 sky130_fd_sc_hd__and4_1 _432_ (.A(_134_),
    .B(net10),
    .C(net42),
    .D(_059_),
    .X(_196_));
 sky130_fd_sc_hd__o2bb2a_4 _433_ (.A1_N(_058_),
    .A2_N(_136_),
    .B1(_196_),
    .B2(_140_),
    .X(\bit_adder[18].FA.sum ));
 sky130_fd_sc_hd__and3_1 _434_ (.A(net43),
    .B(net11),
    .C(_139_),
    .X(_197_));
 sky130_fd_sc_hd__o22a_1 _435_ (.A1(_056_),
    .A2(_139_),
    .B1(_143_),
    .B2(_197_),
    .X(\bit_adder[19].FA.sum ));
 sky130_fd_sc_hd__xnor2_1 _436_ (.A(net45),
    .B(net13),
    .Y(_198_));
 sky130_fd_sc_hd__xor2_1 _437_ (.A(_143_),
    .B(_198_),
    .X(\bit_adder[20].FA.sum ));
 sky130_fd_sc_hd__a21oi_1 _438_ (.A1(_054_),
    .A2(_055_),
    .B1(_146_),
    .Y(_199_));
 sky130_fd_sc_hd__and3_1 _439_ (.A(_146_),
    .B(_055_),
    .C(_054_),
    .X(_200_));
 sky130_fd_sc_hd__nor2_1 _440_ (.A(_199_),
    .B(_200_),
    .Y(\bit_adder[21].FA.sum ));
 sky130_fd_sc_hd__and3_1 _441_ (.A(net47),
    .B(net15),
    .C(_149_),
    .X(_201_));
 sky130_fd_sc_hd__o22a_1 _442_ (.A1(_052_),
    .A2(_149_),
    .B1(_201_),
    .B2(_152_),
    .X(\bit_adder[22].FA.sum ));
 sky130_fd_sc_hd__or3b_1 _443_ (.A(net48),
    .B(net16),
    .C_N(_152_),
    .X(_202_));
 sky130_fd_sc_hd__a2bb2o_1 _444_ (.A1_N(_051_),
    .A2_N(_152_),
    .B1(_155_),
    .B2(_202_),
    .X(\bit_adder[23].FA.sum ));
 sky130_fd_sc_hd__and2_1 _445_ (.A(_049_),
    .B(_050_),
    .X(_203_));
 sky130_fd_sc_hd__xnor2_1 _446_ (.A(_155_),
    .B(_203_),
    .Y(\bit_adder[24].FA.sum ));
 sky130_fd_sc_hd__nand2_1 _447_ (.A(_047_),
    .B(_048_),
    .Y(_204_));
 sky130_fd_sc_hd__xor2_1 _448_ (.A(_158_),
    .B(_204_),
    .X(\bit_adder[25].FA.sum ));
 sky130_fd_sc_hd__a22oi_1 _449_ (.A1(_045_),
    .A2(_046_),
    .B1(_047_),
    .B2(_159_),
    .Y(_205_));
 sky130_fd_sc_hd__and4_1 _450_ (.A(_045_),
    .B(_046_),
    .C(_047_),
    .D(_159_),
    .X(_206_));
 sky130_fd_sc_hd__nor2_1 _451_ (.A(_205_),
    .B(_206_),
    .Y(\bit_adder[26].FA.sum ));
 sky130_fd_sc_hd__and3_1 _452_ (.A(net52),
    .B(net20),
    .C(_163_),
    .X(_207_));
 sky130_fd_sc_hd__o22a_1 _453_ (.A1(_043_),
    .A2(_163_),
    .B1(_166_),
    .B2(_207_),
    .X(\bit_adder[27].FA.sum ));
 sky130_fd_sc_hd__a21oi_1 _454_ (.A1(_041_),
    .A2(_042_),
    .B1(_166_),
    .Y(_208_));
 sky130_fd_sc_hd__and3_1 _455_ (.A(_041_),
    .B(_042_),
    .C(_166_),
    .X(_209_));
 sky130_fd_sc_hd__or2_1 _456_ (.A(_208_),
    .B(_209_),
    .X(\bit_adder[28].FA.sum ));
 sky130_fd_sc_hd__a22oi_1 _457_ (.A1(_039_),
    .A2(_040_),
    .B1(_041_),
    .B2(_167_),
    .Y(_210_));
 sky130_fd_sc_hd__and4_1 _458_ (.A(_039_),
    .B(_040_),
    .C(_041_),
    .D(_167_),
    .X(_211_));
 sky130_fd_sc_hd__nor2_1 _459_ (.A(_210_),
    .B(_211_),
    .Y(\bit_adder[29].FA.sum ));
 sky130_fd_sc_hd__a22o_1 _460_ (.A1(_036_),
    .A2(_038_),
    .B1(_040_),
    .B2(_170_),
    .X(_212_));
 sky130_fd_sc_hd__nand4_1 _461_ (.A(_036_),
    .B(_038_),
    .C(_040_),
    .D(_170_),
    .Y(_213_));
 sky130_fd_sc_hd__nand2_1 _462_ (.A(_212_),
    .B(_213_),
    .Y(\bit_adder[30].FA.sum ));
 sky130_fd_sc_hd__o221ai_1 _463_ (.A1(net56),
    .A2(net24),
    .B1(_032_),
    .B2(_034_),
    .C1(_171_),
    .Y(_214_));
 sky130_fd_sc_hd__o2111ai_1 _464_ (.A1(_000_),
    .A2(_001_),
    .B1(_033_),
    .C1(_035_),
    .D1(_173_),
    .Y(_215_));
 sky130_fd_sc_hd__nand2_1 _465_ (.A(_214_),
    .B(_215_),
    .Y(\bit_adder[31].FA.sum ));
 sky130_fd_sc_hd__buf_1 _466_ (.A(\bit_adder[18].FA.sum ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 _467_ (.A(\bit_adder[19].FA.sum ),
    .X(net78));
 sky130_fd_sc_hd__buf_1 _468_ (.A(\bit_adder[20].FA.sum ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 _469_ (.A(\bit_adder[21].FA.sum ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 _470_ (.A(\bit_adder[22].FA.sum ),
    .X(net82));
 sky130_fd_sc_hd__buf_1 _471_ (.A(\bit_adder[23].FA.sum ),
    .X(net83));
 sky130_fd_sc_hd__buf_1 _472_ (.A(\bit_adder[24].FA.sum ),
    .X(net84));
 sky130_fd_sc_hd__buf_1 _473_ (.A(\bit_adder[25].FA.sum ),
    .X(net85));
 sky130_fd_sc_hd__buf_1 _474_ (.A(\bit_adder[26].FA.sum ),
    .X(net86));
 sky130_fd_sc_hd__buf_1 _475_ (.A(\bit_adder[27].FA.sum ),
    .X(net87));
 sky130_fd_sc_hd__buf_1 _476_ (.A(\bit_adder[28].FA.sum ),
    .X(net88));
 sky130_fd_sc_hd__buf_1 _477_ (.A(\bit_adder[29].FA.sum ),
    .X(net89));
 sky130_fd_sc_hd__buf_1 _478_ (.A(\bit_adder[30].FA.sum ),
    .X(net91));
 sky130_fd_sc_hd__buf_1 _479_ (.A(\bit_adder[31].FA.sum ),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 _480_ (.A(\bit_adder[0].FA.sum ),
    .X(net68));
 sky130_fd_sc_hd__buf_1 _481_ (.A(\bit_adder[1].FA.sum ),
    .X(net79));
 sky130_fd_sc_hd__buf_1 _482_ (.A(\bit_adder[2].FA.sum ),
    .X(net90));
 sky130_fd_sc_hd__buf_1 _483_ (.A(\bit_adder[3].FA.sum ),
    .X(net93));
 sky130_fd_sc_hd__buf_1 _484_ (.A(\bit_adder[4].FA.sum ),
    .X(net94));
 sky130_fd_sc_hd__buf_1 _485_ (.A(\bit_adder[5].FA.sum ),
    .X(net95));
 sky130_fd_sc_hd__buf_1 _486_ (.A(\bit_adder[6].FA.sum ),
    .X(net96));
 sky130_fd_sc_hd__buf_1 _487_ (.A(\bit_adder[7].FA.sum ),
    .X(net97));
 sky130_fd_sc_hd__buf_1 _488_ (.A(\bit_adder[8].FA.sum ),
    .X(net98));
 sky130_fd_sc_hd__buf_1 _489_ (.A(\bit_adder[9].FA.sum ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 _490_ (.A(\bit_adder[10].FA.sum ),
    .X(net69));
 sky130_fd_sc_hd__buf_1 _491_ (.A(\bit_adder[11].FA.sum ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 _492_ (.A(\bit_adder[12].FA.sum ),
    .X(net71));
 sky130_fd_sc_hd__buf_1 _493_ (.A(\bit_adder[13].FA.sum ),
    .X(net72));
 sky130_fd_sc_hd__buf_1 _494_ (.A(\bit_adder[14].FA.sum ),
    .X(net73));
 sky130_fd_sc_hd__buf_1 _495_ (.A(\bit_adder[15].FA.sum ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 _496_ (.A(\bit_adder[16].FA.sum ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 _497_ (.A(\bit_adder[17].FA.sum ),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(b[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(b[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(b[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_2 input36 (.A(b[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(b[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(b[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(b[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input40 (.A(b[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_4 input41 (.A(b[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(b[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(b[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(b[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(b[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(b[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(b[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(b[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(b[24]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(b[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(b[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(b[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(b[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(b[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(b[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(b[30]),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(b[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(b[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(b[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input60 (.A(b[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 input61 (.A(b[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(b[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(b[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(b[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(cin),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_16 output66 (.A(net66),
    .X(cout));
 sky130_fd_sc_hd__clkbuf_16 output67 (.A(net67),
    .X(overflow));
 sky130_fd_sc_hd__clkbuf_16 output68 (.A(net68),
    .X(sum[0]));
 sky130_fd_sc_hd__clkbuf_16 output69 (.A(net69),
    .X(sum[10]));
 sky130_fd_sc_hd__clkbuf_16 output70 (.A(net70),
    .X(sum[11]));
 sky130_fd_sc_hd__clkbuf_16 output71 (.A(net71),
    .X(sum[12]));
 sky130_fd_sc_hd__clkbuf_16 output72 (.A(net72),
    .X(sum[13]));
 sky130_fd_sc_hd__clkbuf_16 output73 (.A(net73),
    .X(sum[14]));
 sky130_fd_sc_hd__clkbuf_16 output74 (.A(net74),
    .X(sum[15]));
 sky130_fd_sc_hd__clkbuf_16 output75 (.A(net75),
    .X(sum[16]));
 sky130_fd_sc_hd__clkbuf_16 output76 (.A(net76),
    .X(sum[17]));
 sky130_fd_sc_hd__clkbuf_16 output77 (.A(net77),
    .X(sum[18]));
 sky130_fd_sc_hd__clkbuf_16 output78 (.A(net78),
    .X(sum[19]));
 sky130_fd_sc_hd__clkbuf_16 output79 (.A(net79),
    .X(sum[1]));
 sky130_fd_sc_hd__clkbuf_16 output80 (.A(net80),
    .X(sum[20]));
 sky130_fd_sc_hd__clkbuf_16 output81 (.A(net81),
    .X(sum[21]));
 sky130_fd_sc_hd__clkbuf_16 output82 (.A(net82),
    .X(sum[22]));
 sky130_fd_sc_hd__clkbuf_16 output83 (.A(net83),
    .X(sum[23]));
 sky130_fd_sc_hd__clkbuf_16 output84 (.A(net84),
    .X(sum[24]));
 sky130_fd_sc_hd__clkbuf_16 output85 (.A(net85),
    .X(sum[25]));
 sky130_fd_sc_hd__clkbuf_16 output86 (.A(net86),
    .X(sum[26]));
 sky130_fd_sc_hd__clkbuf_16 output87 (.A(net87),
    .X(sum[27]));
 sky130_fd_sc_hd__clkbuf_16 output88 (.A(net88),
    .X(sum[28]));
 sky130_fd_sc_hd__clkbuf_16 output89 (.A(net89),
    .X(sum[29]));
 sky130_fd_sc_hd__clkbuf_16 output90 (.A(net90),
    .X(sum[2]));
 sky130_fd_sc_hd__clkbuf_16 output91 (.A(net91),
    .X(sum[30]));
 sky130_fd_sc_hd__clkbuf_16 output92 (.A(net92),
    .X(sum[31]));
 sky130_fd_sc_hd__clkbuf_16 output93 (.A(net93),
    .X(sum[3]));
 sky130_fd_sc_hd__clkbuf_16 output94 (.A(net94),
    .X(sum[4]));
 sky130_fd_sc_hd__clkbuf_16 output95 (.A(net95),
    .X(sum[5]));
 sky130_fd_sc_hd__clkbuf_16 output96 (.A(net96),
    .X(sum[6]));
 sky130_fd_sc_hd__clkbuf_16 output97 (.A(net97),
    .X(sum[7]));
 sky130_fd_sc_hd__clkbuf_16 output98 (.A(net98),
    .X(sum[8]));
 sky130_fd_sc_hd__clkbuf_16 output99 (.A(net99),
    .X(sum[9]));
endmodule
