module carry_bypass_adder_routing(cin,
    clk,
    cout,
    overflow,
    a,
    b,
    sum);
 input cin;
 input clk;
 output cout;
 output overflow;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire \carry_ripple[0].RA.full_adder[0].FA.out ;
 wire \carry_ripple[0].RA.full_adder[1].FA.out ;
 wire \carry_ripple[0].RA.full_adder[2].FA.out ;
 wire \carry_ripple[0].RA.full_adder[3].FA.out ;
 wire \carry_ripple[1].RA.full_adder[0].FA.out ;
 wire \carry_ripple[1].RA.full_adder[1].FA.out ;
 wire \carry_ripple[1].RA.full_adder[2].FA.out ;
 wire \carry_ripple[1].RA.full_adder[3].FA.out ;
 wire \carry_ripple[2].RA.full_adder[0].FA.out ;
 wire \carry_ripple[2].RA.full_adder[1].FA.out ;
 wire \carry_ripple[2].RA.full_adder[2].FA.out ;
 wire \carry_ripple[2].RA.full_adder[3].FA.out ;
 wire \carry_ripple[3].RA.full_adder[0].FA.out ;
 wire \carry_ripple[3].RA.full_adder[1].FA.out ;
 wire \carry_ripple[3].RA.full_adder[2].FA.out ;
 wire \carry_ripple[3].RA.full_adder[3].FA.out ;
 wire \carry_ripple[4].RA.full_adder[0].FA.out ;
 wire \carry_ripple[4].RA.full_adder[1].FA.out ;
 wire \carry_ripple[4].RA.full_adder[2].FA.out ;
 wire \carry_ripple[4].RA.full_adder[3].FA.out ;
 wire \carry_ripple[5].RA.full_adder[0].FA.out ;
 wire \carry_ripple[5].RA.full_adder[1].FA.out ;
 wire \carry_ripple[5].RA.full_adder[2].FA.out ;
 wire \carry_ripple[5].RA.full_adder[3].FA.out ;
 wire \carry_ripple[6].RA.full_adder[0].FA.out ;
 wire \carry_ripple[6].RA.full_adder[1].FA.out ;
 wire \carry_ripple[6].RA.full_adder[2].FA.out ;
 wire \carry_ripple[6].RA.full_adder[3].FA.out ;
 wire \carry_ripple[7].RA.full_adder[0].FA.out ;
 wire \carry_ripple[7].RA.full_adder[1].FA.out ;
 wire \carry_ripple[7].RA.full_adder[2].FA.out ;
 wire \carry_ripple[7].RA.full_adder[3].FA.out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__inv_2 _194_ (.A(net56),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _195_ (.A(net24),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _196_ (.A(net58),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _197_ (.A(net26),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _198_ (.A(net44),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _199_ (.A(net12),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _200_ (.A(net60),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _201_ (.A(net28),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _202_ (.A(net64),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _203_ (.A(net32),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _204_ (.A(net63),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _205_ (.A(net31),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _206_ (.A(net37),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _207_ (.A(net5),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _208_ (.A(net41),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _209_ (.A(net9),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _210_ (.A(net46),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _211_ (.A(net14),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _212_ (.A(net50),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _213_ (.A(net18),
    .Y(_019_));
 sky130_fd_sc_hd__nor2_1 _214_ (.A(net57),
    .B(net25),
    .Y(_020_));
 sky130_fd_sc_hd__and2_1 _215_ (.A(net57),
    .B(net25),
    .X(_021_));
 sky130_fd_sc_hd__nand2_1 _216_ (.A(net57),
    .B(net25),
    .Y(_022_));
 sky130_fd_sc_hd__nor2_1 _217_ (.A(_020_),
    .B(_021_),
    .Y(_023_));
 sky130_fd_sc_hd__nor2_1 _218_ (.A(_000_),
    .B(_001_),
    .Y(_024_));
 sky130_fd_sc_hd__nor2_1 _219_ (.A(net56),
    .B(net24),
    .Y(_025_));
 sky130_fd_sc_hd__or2_1 _220_ (.A(net56),
    .B(net24),
    .X(_026_));
 sky130_fd_sc_hd__and2_1 _221_ (.A(net54),
    .B(net22),
    .X(_027_));
 sky130_fd_sc_hd__nand2_2 _222_ (.A(net54),
    .B(net22),
    .Y(_028_));
 sky130_fd_sc_hd__or2_1 _223_ (.A(net54),
    .B(net22),
    .X(_029_));
 sky130_fd_sc_hd__and2_2 _224_ (.A(net53),
    .B(net21),
    .X(_030_));
 sky130_fd_sc_hd__nor2_1 _225_ (.A(net53),
    .B(net21),
    .Y(_031_));
 sky130_fd_sc_hd__or2_1 _226_ (.A(net53),
    .B(net21),
    .X(_032_));
 sky130_fd_sc_hd__nor2_1 _227_ (.A(net49),
    .B(net17),
    .Y(_033_));
 sky130_fd_sc_hd__and2_1 _228_ (.A(net49),
    .B(net17),
    .X(_034_));
 sky130_fd_sc_hd__nor2_1 _229_ (.A(_033_),
    .B(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__or2_1 _230_ (.A(net51),
    .B(net19),
    .X(_036_));
 sky130_fd_sc_hd__nand2_1 _231_ (.A(net51),
    .B(net19),
    .Y(_037_));
 sky130_fd_sc_hd__and2_1 _232_ (.A(_036_),
    .B(_037_),
    .X(_038_));
 sky130_fd_sc_hd__xor2_1 _233_ (.A(net50),
    .B(net18),
    .X(_039_));
 sky130_fd_sc_hd__xor2_1 _234_ (.A(net52),
    .B(net20),
    .X(_040_));
 sky130_fd_sc_hd__nand4_1 _235_ (.A(_035_),
    .B(_038_),
    .C(_039_),
    .D(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _236_ (.A(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__nor2_2 _237_ (.A(net45),
    .B(net13),
    .Y(_043_));
 sky130_fd_sc_hd__and2_2 _238_ (.A(net45),
    .B(net13),
    .X(_044_));
 sky130_fd_sc_hd__nor2_1 _239_ (.A(_043_),
    .B(_044_),
    .Y(_045_));
 sky130_fd_sc_hd__or2_1 _240_ (.A(net47),
    .B(net15),
    .X(_046_));
 sky130_fd_sc_hd__nand2_1 _241_ (.A(net47),
    .B(net15),
    .Y(_047_));
 sky130_fd_sc_hd__and2_1 _242_ (.A(_046_),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__xor2_4 _243_ (.A(net46),
    .B(net14),
    .X(_049_));
 sky130_fd_sc_hd__xor2_1 _244_ (.A(net48),
    .B(net16),
    .X(_050_));
 sky130_fd_sc_hd__nand4_1 _245_ (.A(_045_),
    .B(_048_),
    .C(_049_),
    .D(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _246_ (.A(_051_),
    .Y(_052_));
 sky130_fd_sc_hd__nor2_1 _247_ (.A(net40),
    .B(net8),
    .Y(_053_));
 sky130_fd_sc_hd__and2_1 _248_ (.A(net40),
    .B(net8),
    .X(_054_));
 sky130_fd_sc_hd__nor2_1 _249_ (.A(_053_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__or2_1 _250_ (.A(net42),
    .B(net10),
    .X(_056_));
 sky130_fd_sc_hd__nand2_1 _251_ (.A(net42),
    .B(net10),
    .Y(_057_));
 sky130_fd_sc_hd__and2_1 _252_ (.A(_056_),
    .B(_057_),
    .X(_058_));
 sky130_fd_sc_hd__xor2_2 _253_ (.A(net41),
    .B(net9),
    .X(_059_));
 sky130_fd_sc_hd__xor2_4 _254_ (.A(net43),
    .B(net11),
    .X(_060_));
 sky130_fd_sc_hd__and4_4 _255_ (.A(_055_),
    .B(_058_),
    .C(_059_),
    .D(_060_),
    .X(_061_));
 sky130_fd_sc_hd__or2_2 _256_ (.A(net38),
    .B(net6),
    .X(_062_));
 sky130_fd_sc_hd__nand2_1 _257_ (.A(net38),
    .B(net6),
    .Y(_063_));
 sky130_fd_sc_hd__and2_4 _258_ (.A(net36),
    .B(net4),
    .X(_064_));
 sky130_fd_sc_hd__or2_1 _259_ (.A(net61),
    .B(net29),
    .X(_065_));
 sky130_fd_sc_hd__nand2_1 _260_ (.A(net61),
    .B(net29),
    .Y(_066_));
 sky130_fd_sc_hd__and2_1 _261_ (.A(_065_),
    .B(_066_),
    .X(_067_));
 sky130_fd_sc_hd__or2_1 _262_ (.A(net59),
    .B(net27),
    .X(_068_));
 sky130_fd_sc_hd__nand2_1 _263_ (.A(net59),
    .B(net27),
    .Y(_069_));
 sky130_fd_sc_hd__and2_1 _264_ (.A(_068_),
    .B(_069_),
    .X(_070_));
 sky130_fd_sc_hd__xor2_1 _265_ (.A(net62),
    .B(net30),
    .X(_071_));
 sky130_fd_sc_hd__nor2_1 _266_ (.A(net60),
    .B(net28),
    .Y(_072_));
 sky130_fd_sc_hd__nor2_1 _267_ (.A(_006_),
    .B(_007_),
    .Y(_073_));
 sky130_fd_sc_hd__nor2_1 _268_ (.A(_072_),
    .B(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__nand4_1 _269_ (.A(_067_),
    .B(_070_),
    .C(_071_),
    .D(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _270_ (.A(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__or2_1 _271_ (.A(net58),
    .B(net26),
    .X(_077_));
 sky130_fd_sc_hd__nand2_1 _272_ (.A(net58),
    .B(net26),
    .Y(_078_));
 sky130_fd_sc_hd__nor2_1 _273_ (.A(net55),
    .B(net23),
    .Y(_079_));
 sky130_fd_sc_hd__nand2_1 _274_ (.A(net55),
    .B(net23),
    .Y(_080_));
 sky130_fd_sc_hd__or2_1 _275_ (.A(net33),
    .B(net1),
    .X(_081_));
 sky130_fd_sc_hd__a21o_1 _276_ (.A1(net33),
    .A2(net1),
    .B1(net65),
    .X(_082_));
 sky130_fd_sc_hd__o21a_1 _277_ (.A1(net33),
    .A2(net1),
    .B1(net65),
    .X(_083_));
 sky130_fd_sc_hd__o21ai_1 _278_ (.A1(net33),
    .A2(net1),
    .B1(_082_),
    .Y(_084_));
 sky130_fd_sc_hd__a221o_1 _279_ (.A1(net44),
    .A2(net12),
    .B1(net33),
    .B2(net1),
    .C1(_083_),
    .X(_085_));
 sky130_fd_sc_hd__o221ai_4 _280_ (.A1(net44),
    .A2(net12),
    .B1(net33),
    .B2(net1),
    .C1(_082_),
    .Y(_086_));
 sky130_fd_sc_hd__o21a_1 _281_ (.A1(_004_),
    .A2(_005_),
    .B1(_086_),
    .X(_087_));
 sky130_fd_sc_hd__o211ai_2 _282_ (.A1(_004_),
    .A2(_005_),
    .B1(_080_),
    .C1(_086_),
    .Y(_088_));
 sky130_fd_sc_hd__o21ai_1 _283_ (.A1(net55),
    .A2(net23),
    .B1(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__o211ai_2 _284_ (.A1(net55),
    .A2(net23),
    .B1(_077_),
    .C1(_088_),
    .Y(_090_));
 sky130_fd_sc_hd__o21a_1 _285_ (.A1(_002_),
    .A2(_003_),
    .B1(_090_),
    .X(_091_));
 sky130_fd_sc_hd__nand2_1 _286_ (.A(_076_),
    .B(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__o211ai_2 _287_ (.A1(_002_),
    .A2(_003_),
    .B1(_069_),
    .C1(_090_),
    .Y(_093_));
 sky130_fd_sc_hd__o211ai_1 _288_ (.A1(net60),
    .A2(net28),
    .B1(_068_),
    .C1(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__a22o_1 _289_ (.A1(net60),
    .A2(net28),
    .B1(_068_),
    .B2(_093_),
    .X(_095_));
 sky130_fd_sc_hd__o21a_1 _290_ (.A1(_006_),
    .A2(_007_),
    .B1(_094_),
    .X(_096_));
 sky130_fd_sc_hd__o211ai_1 _291_ (.A1(_006_),
    .A2(_007_),
    .B1(_066_),
    .C1(_094_),
    .Y(_097_));
 sky130_fd_sc_hd__o21ai_1 _292_ (.A1(net61),
    .A2(net29),
    .B1(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__o211ai_1 _293_ (.A1(net62),
    .A2(net30),
    .B1(_065_),
    .C1(_097_),
    .Y(_099_));
 sky130_fd_sc_hd__a21oi_1 _294_ (.A1(net62),
    .A2(net30),
    .B1(_076_),
    .Y(_100_));
 sky130_fd_sc_hd__nand2_1 _295_ (.A(_099_),
    .B(_100_),
    .Y(_101_));
 sky130_fd_sc_hd__a22o_2 _296_ (.A1(_076_),
    .A2(_091_),
    .B1(_099_),
    .B2(_100_),
    .X(_102_));
 sky130_fd_sc_hd__xor2_1 _297_ (.A(net63),
    .B(net31),
    .X(_103_));
 sky130_fd_sc_hd__or2_1 _298_ (.A(net34),
    .B(net2),
    .X(_104_));
 sky130_fd_sc_hd__nand2_1 _299_ (.A(net34),
    .B(net2),
    .Y(_105_));
 sky130_fd_sc_hd__and2_1 _300_ (.A(_104_),
    .B(_105_),
    .X(_106_));
 sky130_fd_sc_hd__xor2_2 _301_ (.A(net64),
    .B(net32),
    .X(_107_));
 sky130_fd_sc_hd__xor2_1 _302_ (.A(net35),
    .B(net3),
    .X(_108_));
 sky130_fd_sc_hd__nand4_1 _303_ (.A(_103_),
    .B(_106_),
    .C(_107_),
    .D(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _304_ (.A(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__a2bb2oi_2 _305_ (.A1_N(_010_),
    .A2_N(_011_),
    .B1(_092_),
    .B2(_101_),
    .Y(_111_));
 sky130_fd_sc_hd__a22o_1 _306_ (.A1(_008_),
    .A2(_009_),
    .B1(_010_),
    .B2(_011_),
    .X(_112_));
 sky130_fd_sc_hd__o22a_1 _307_ (.A1(_008_),
    .A2(_009_),
    .B1(_112_),
    .B2(_111_),
    .X(_113_));
 sky130_fd_sc_hd__o221ai_4 _308_ (.A1(_008_),
    .A2(_009_),
    .B1(_112_),
    .B2(_111_),
    .C1(_105_),
    .Y(_114_));
 sky130_fd_sc_hd__o21ai_1 _309_ (.A1(net34),
    .A2(net2),
    .B1(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__o211ai_4 _310_ (.A1(net35),
    .A2(net3),
    .B1(_104_),
    .C1(_114_),
    .Y(_116_));
 sky130_fd_sc_hd__a21oi_2 _311_ (.A1(net35),
    .A2(net3),
    .B1(_110_),
    .Y(_117_));
 sky130_fd_sc_hd__a22oi_4 _312_ (.A1(_102_),
    .A2(_110_),
    .B1(_116_),
    .B2(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__a22o_4 _313_ (.A1(_102_),
    .A2(_110_),
    .B1(_116_),
    .B2(_117_),
    .X(_119_));
 sky130_fd_sc_hd__a21o_1 _314_ (.A1(net36),
    .A2(net4),
    .B1(_118_),
    .X(_120_));
 sky130_fd_sc_hd__nor2_4 _315_ (.A(net36),
    .B(net4),
    .Y(_121_));
 sky130_fd_sc_hd__a21o_1 _316_ (.A1(_012_),
    .A2(_013_),
    .B1(_121_),
    .X(_122_));
 sky130_fd_sc_hd__o21bai_2 _317_ (.A1(_064_),
    .A2(_118_),
    .B1_N(_122_),
    .Y(_123_));
 sky130_fd_sc_hd__o21a_1 _318_ (.A1(_012_),
    .A2(_013_),
    .B1(_123_),
    .X(_124_));
 sky130_fd_sc_hd__o211ai_4 _319_ (.A1(_012_),
    .A2(_013_),
    .B1(_063_),
    .C1(_123_),
    .Y(_125_));
 sky130_fd_sc_hd__o211ai_4 _320_ (.A1(net39),
    .A2(net7),
    .B1(_062_),
    .C1(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__xor2_1 _321_ (.A(net37),
    .B(net5),
    .X(_127_));
 sky130_fd_sc_hd__nor2_4 _322_ (.A(_064_),
    .B(_121_),
    .Y(_128_));
 sky130_fd_sc_hd__xor2_1 _323_ (.A(net39),
    .B(net7),
    .X(_129_));
 sky130_fd_sc_hd__and2_1 _324_ (.A(_062_),
    .B(_063_),
    .X(_130_));
 sky130_fd_sc_hd__nand4_1 _325_ (.A(_127_),
    .B(_128_),
    .C(_129_),
    .D(_130_),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _326_ (.A(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__a21oi_2 _327_ (.A1(net39),
    .A2(net7),
    .B1(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__a22oi_4 _328_ (.A1(_119_),
    .A2(_132_),
    .B1(_126_),
    .B2(_133_),
    .Y(_134_));
 sky130_fd_sc_hd__a22o_4 _329_ (.A1(_119_),
    .A2(_132_),
    .B1(_126_),
    .B2(_133_),
    .X(_135_));
 sky130_fd_sc_hd__a21o_1 _330_ (.A1(_014_),
    .A2(_015_),
    .B1(_053_),
    .X(_136_));
 sky130_fd_sc_hd__o21bai_2 _331_ (.A1(_054_),
    .A2(_134_),
    .B1_N(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__o21a_1 _332_ (.A1(_014_),
    .A2(_015_),
    .B1(_137_),
    .X(_138_));
 sky130_fd_sc_hd__o211ai_4 _333_ (.A1(_014_),
    .A2(_015_),
    .B1(_057_),
    .C1(_137_),
    .Y(_139_));
 sky130_fd_sc_hd__o21ai_2 _334_ (.A1(net42),
    .A2(net10),
    .B1(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__o211ai_4 _335_ (.A1(net43),
    .A2(net11),
    .B1(_056_),
    .C1(_139_),
    .Y(_141_));
 sky130_fd_sc_hd__a21oi_2 _336_ (.A1(net43),
    .A2(net11),
    .B1(_061_),
    .Y(_142_));
 sky130_fd_sc_hd__a22oi_4 _337_ (.A1(_061_),
    .A2(_135_),
    .B1(_141_),
    .B2(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__a22o_2 _338_ (.A1(_061_),
    .A2(_135_),
    .B1(_141_),
    .B2(_142_),
    .X(_144_));
 sky130_fd_sc_hd__a21o_1 _339_ (.A1(_016_),
    .A2(_017_),
    .B1(_043_),
    .X(_145_));
 sky130_fd_sc_hd__o21bai_1 _340_ (.A1(_044_),
    .A2(_143_),
    .B1_N(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__o21ai_1 _341_ (.A1(_016_),
    .A2(_017_),
    .B1(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__o211ai_2 _342_ (.A1(_016_),
    .A2(_017_),
    .B1(_047_),
    .C1(_146_),
    .Y(_148_));
 sky130_fd_sc_hd__o21ai_1 _343_ (.A1(net47),
    .A2(net15),
    .B1(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__o211ai_4 _344_ (.A1(net48),
    .A2(net16),
    .B1(_046_),
    .C1(_148_),
    .Y(_150_));
 sky130_fd_sc_hd__a21oi_2 _345_ (.A1(net48),
    .A2(net16),
    .B1(_052_),
    .Y(_151_));
 sky130_fd_sc_hd__a22oi_4 _346_ (.A1(_052_),
    .A2(_144_),
    .B1(_150_),
    .B2(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__a22o_2 _347_ (.A1(_052_),
    .A2(_144_),
    .B1(_150_),
    .B2(_151_),
    .X(_153_));
 sky130_fd_sc_hd__a21oi_1 _348_ (.A1(net49),
    .A2(net17),
    .B1(_152_),
    .Y(_154_));
 sky130_fd_sc_hd__a21o_1 _349_ (.A1(_018_),
    .A2(_019_),
    .B1(_033_),
    .X(_155_));
 sky130_fd_sc_hd__o21bai_1 _350_ (.A1(_034_),
    .A2(_152_),
    .B1_N(_155_),
    .Y(_156_));
 sky130_fd_sc_hd__o22a_1 _351_ (.A1(_018_),
    .A2(_019_),
    .B1(_155_),
    .B2(_154_),
    .X(_157_));
 sky130_fd_sc_hd__o211ai_2 _352_ (.A1(_018_),
    .A2(_019_),
    .B1(_037_),
    .C1(_156_),
    .Y(_158_));
 sky130_fd_sc_hd__o21ai_1 _353_ (.A1(net51),
    .A2(net19),
    .B1(_158_),
    .Y(_159_));
 sky130_fd_sc_hd__o211ai_4 _354_ (.A1(net52),
    .A2(net20),
    .B1(_036_),
    .C1(_158_),
    .Y(_160_));
 sky130_fd_sc_hd__a21oi_2 _355_ (.A1(net52),
    .A2(net20),
    .B1(_042_),
    .Y(_161_));
 sky130_fd_sc_hd__a22oi_4 _356_ (.A1(_042_),
    .A2(_153_),
    .B1(_160_),
    .B2(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__a221oi_2 _357_ (.A1(_042_),
    .A2(_153_),
    .B1(_160_),
    .B2(_161_),
    .C1(_031_),
    .Y(_163_));
 sky130_fd_sc_hd__o21ai_1 _358_ (.A1(_030_),
    .A2(_162_),
    .B1(_032_),
    .Y(_164_));
 sky130_fd_sc_hd__o221ai_4 _359_ (.A1(net54),
    .A2(net22),
    .B1(_030_),
    .B2(_162_),
    .C1(_032_),
    .Y(_165_));
 sky130_fd_sc_hd__a2bb2oi_1 _360_ (.A1_N(net56),
    .A2_N(net24),
    .B1(_028_),
    .B2(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__o311ai_2 _361_ (.A1(_027_),
    .A2(_030_),
    .A3(_163_),
    .B1(_029_),
    .C1(_026_),
    .Y(_167_));
 sky130_fd_sc_hd__o211ai_4 _362_ (.A1(_000_),
    .A2(_001_),
    .B1(_028_),
    .C1(_165_),
    .Y(_168_));
 sky130_fd_sc_hd__o21ai_1 _363_ (.A1(net56),
    .A2(net24),
    .B1(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__o221ai_1 _364_ (.A1(net56),
    .A2(net24),
    .B1(_020_),
    .B2(_021_),
    .C1(_168_),
    .Y(_170_));
 sky130_fd_sc_hd__o211ai_1 _365_ (.A1(_000_),
    .A2(_001_),
    .B1(_023_),
    .C1(_167_),
    .Y(_171_));
 sky130_fd_sc_hd__nand2_1 _366_ (.A(_170_),
    .B(_171_),
    .Y(\carry_ripple[7].RA.full_adder[3].FA.out ));
 sky130_fd_sc_hd__o221ai_1 _367_ (.A1(net57),
    .A2(net25),
    .B1(net56),
    .B2(net24),
    .C1(_168_),
    .Y(_172_));
 sky130_fd_sc_hd__o31a_1 _368_ (.A1(_021_),
    .A2(_024_),
    .A3(_166_),
    .B1(_172_),
    .X(net67));
 sky130_fd_sc_hd__nor2_1 _369_ (.A(_030_),
    .B(_031_),
    .Y(_173_));
 sky130_fd_sc_hd__nand2_1 _370_ (.A(_028_),
    .B(_029_),
    .Y(_174_));
 sky130_fd_sc_hd__or4_1 _371_ (.A(_024_),
    .B(_025_),
    .C(_030_),
    .D(_031_),
    .X(_175_));
 sky130_fd_sc_hd__or3_1 _372_ (.A(_021_),
    .B(_174_),
    .C(_175_),
    .X(_176_));
 sky130_fd_sc_hd__o22ai_1 _373_ (.A1(net57),
    .A2(net25),
    .B1(_176_),
    .B2(_162_),
    .Y(_177_));
 sky130_fd_sc_hd__a31oi_2 _374_ (.A1(_169_),
    .A2(_176_),
    .A3(_022_),
    .B1(_177_),
    .Y(net66));
 sky130_fd_sc_hd__o2111ai_1 _375_ (.A1(_079_),
    .A2(_087_),
    .B1(_080_),
    .C1(_002_),
    .D1(_003_),
    .Y(_178_));
 sky130_fd_sc_hd__a2bb2o_1 _376_ (.A1_N(_078_),
    .A2_N(_089_),
    .B1(_091_),
    .B2(_178_),
    .X(\carry_ripple[0].RA.full_adder[3].FA.out ));
 sky130_fd_sc_hd__o2111a_1 _377_ (.A1(net44),
    .A2(net12),
    .B1(net55),
    .C1(net23),
    .D1(_085_),
    .X(_179_));
 sky130_fd_sc_hd__o2bb2a_1 _378_ (.A1_N(_079_),
    .A2_N(_087_),
    .B1(_089_),
    .B2(_179_),
    .X(\carry_ripple[0].RA.full_adder[2].FA.out ));
 sky130_fd_sc_hd__and4_1 _379_ (.A(_081_),
    .B(_082_),
    .C(net44),
    .D(net12),
    .X(_180_));
 sky130_fd_sc_hd__a2111o_1 _380_ (.A1(net33),
    .A2(net1),
    .B1(_083_),
    .C1(net12),
    .D1(net44),
    .X(_181_));
 sky130_fd_sc_hd__a21o_1 _381_ (.A1(_087_),
    .A2(_181_),
    .B1(_180_),
    .X(\carry_ripple[0].RA.full_adder[1].FA.out ));
 sky130_fd_sc_hd__and3_1 _382_ (.A(net65),
    .B(net33),
    .C(net1),
    .X(_182_));
 sky130_fd_sc_hd__or2_1 _383_ (.A(_182_),
    .B(_084_),
    .X(_183_));
 sky130_fd_sc_hd__o21a_1 _384_ (.A1(net65),
    .A2(_081_),
    .B1(_183_),
    .X(\carry_ripple[0].RA.full_adder[0].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _385_ (.A(_071_),
    .B(_098_),
    .Y(\carry_ripple[1].RA.full_adder[3].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _386_ (.A(_067_),
    .B(_096_),
    .Y(\carry_ripple[1].RA.full_adder[2].FA.out ));
 sky130_fd_sc_hd__o221ai_1 _387_ (.A1(net59),
    .A2(net27),
    .B1(_072_),
    .B2(_073_),
    .C1(_093_),
    .Y(_184_));
 sky130_fd_sc_hd__o21ai_1 _388_ (.A1(_072_),
    .A2(_095_),
    .B1(_184_),
    .Y(\carry_ripple[1].RA.full_adder[1].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _389_ (.A(_070_),
    .B(_091_),
    .Y(\carry_ripple[1].RA.full_adder[0].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _390_ (.A(_108_),
    .B(_115_),
    .Y(\carry_ripple[2].RA.full_adder[3].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _391_ (.A(_106_),
    .B(_113_),
    .Y(\carry_ripple[2].RA.full_adder[2].FA.out ));
 sky130_fd_sc_hd__a21o_1 _392_ (.A1(_010_),
    .A2(_011_),
    .B1(_111_),
    .X(_185_));
 sky130_fd_sc_hd__xnor2_1 _393_ (.A(_107_),
    .B(_185_),
    .Y(\carry_ripple[2].RA.full_adder[1].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _394_ (.A(_102_),
    .B(_103_),
    .Y(\carry_ripple[2].RA.full_adder[0].FA.out ));
 sky130_fd_sc_hd__a21oi_1 _395_ (.A1(_062_),
    .A2(_125_),
    .B1(_129_),
    .Y(_186_));
 sky130_fd_sc_hd__and3_1 _396_ (.A(_062_),
    .B(_125_),
    .C(_129_),
    .X(_187_));
 sky130_fd_sc_hd__nor2_1 _397_ (.A(_186_),
    .B(_187_),
    .Y(\carry_ripple[3].RA.full_adder[3].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _398_ (.A(_124_),
    .B(_130_),
    .Y(\carry_ripple[3].RA.full_adder[2].FA.out ));
 sky130_fd_sc_hd__o21a_4 _399_ (.A1(net36),
    .A2(net4),
    .B1(_120_),
    .X(_188_));
 sky130_fd_sc_hd__xor2_1 _400_ (.A(_127_),
    .B(_188_),
    .X(\carry_ripple[3].RA.full_adder[1].FA.out ));
 sky130_fd_sc_hd__a221o_1 _401_ (.A1(_102_),
    .A2(_110_),
    .B1(_116_),
    .B2(_117_),
    .C1(_128_),
    .X(_189_));
 sky130_fd_sc_hd__o21ai_1 _402_ (.A1(_121_),
    .A2(_120_),
    .B1(_189_),
    .Y(\carry_ripple[3].RA.full_adder[0].FA.out ));
 sky130_fd_sc_hd__xnor2_4 _403_ (.A(_060_),
    .B(_140_),
    .Y(\carry_ripple[4].RA.full_adder[3].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _404_ (.A(_058_),
    .B(_138_),
    .Y(\carry_ripple[4].RA.full_adder[2].FA.out ));
 sky130_fd_sc_hd__o21ba_1 _405_ (.A1(_054_),
    .A2(_134_),
    .B1_N(_053_),
    .X(_190_));
 sky130_fd_sc_hd__xor2_1 _406_ (.A(_059_),
    .B(_190_),
    .X(\carry_ripple[4].RA.full_adder[1].FA.out ));
 sky130_fd_sc_hd__xor2_1 _407_ (.A(_055_),
    .B(_134_),
    .X(\carry_ripple[4].RA.full_adder[0].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _408_ (.A(_050_),
    .B(_149_),
    .Y(\carry_ripple[5].RA.full_adder[3].FA.out ));
 sky130_fd_sc_hd__xor2_1 _409_ (.A(_048_),
    .B(_147_),
    .X(\carry_ripple[5].RA.full_adder[2].FA.out ));
 sky130_fd_sc_hd__o21ba_1 _410_ (.A1(_044_),
    .A2(_143_),
    .B1_N(_043_),
    .X(_191_));
 sky130_fd_sc_hd__xor2_1 _411_ (.A(_049_),
    .B(_191_),
    .X(\carry_ripple[5].RA.full_adder[1].FA.out ));
 sky130_fd_sc_hd__xor2_1 _412_ (.A(_045_),
    .B(_143_),
    .X(\carry_ripple[5].RA.full_adder[0].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _413_ (.A(_040_),
    .B(_159_),
    .Y(\carry_ripple[6].RA.full_adder[3].FA.out ));
 sky130_fd_sc_hd__xnor2_1 _414_ (.A(_038_),
    .B(_157_),
    .Y(\carry_ripple[6].RA.full_adder[2].FA.out ));
 sky130_fd_sc_hd__or2_1 _415_ (.A(_033_),
    .B(_154_),
    .X(_192_));
 sky130_fd_sc_hd__xnor2_1 _416_ (.A(_039_),
    .B(_192_),
    .Y(\carry_ripple[6].RA.full_adder[1].FA.out ));
 sky130_fd_sc_hd__xor2_1 _417_ (.A(_035_),
    .B(_152_),
    .X(\carry_ripple[6].RA.full_adder[0].FA.out ));
 sky130_fd_sc_hd__a2bb2oi_1 _418_ (.A1_N(_024_),
    .A2_N(_025_),
    .B1(_028_),
    .B2(_165_),
    .Y(_193_));
 sky130_fd_sc_hd__o21bai_1 _419_ (.A1(_025_),
    .A2(_168_),
    .B1_N(_193_),
    .Y(\carry_ripple[7].RA.full_adder[2].FA.out ));
 sky130_fd_sc_hd__xor2_1 _420_ (.A(_164_),
    .B(_174_),
    .X(\carry_ripple[7].RA.full_adder[1].FA.out ));
 sky130_fd_sc_hd__xor2_1 _421_ (.A(_162_),
    .B(_173_),
    .X(\carry_ripple[7].RA.full_adder[0].FA.out ));
 sky130_fd_sc_hd__buf_1 _422_ (.A(\carry_ripple[0].RA.full_adder[0].FA.out ),
    .X(net68));
 sky130_fd_sc_hd__buf_1 _423_ (.A(\carry_ripple[0].RA.full_adder[1].FA.out ),
    .X(net79));
 sky130_fd_sc_hd__buf_1 _424_ (.A(\carry_ripple[0].RA.full_adder[2].FA.out ),
    .X(net90));
 sky130_fd_sc_hd__buf_1 _425_ (.A(\carry_ripple[0].RA.full_adder[3].FA.out ),
    .X(net93));
 sky130_fd_sc_hd__buf_1 _426_ (.A(\carry_ripple[1].RA.full_adder[0].FA.out ),
    .X(net94));
 sky130_fd_sc_hd__buf_1 _427_ (.A(\carry_ripple[1].RA.full_adder[1].FA.out ),
    .X(net95));
 sky130_fd_sc_hd__buf_1 _428_ (.A(\carry_ripple[1].RA.full_adder[2].FA.out ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _429_ (.A(\carry_ripple[1].RA.full_adder[3].FA.out ),
    .X(net97));
 sky130_fd_sc_hd__buf_1 _430_ (.A(\carry_ripple[2].RA.full_adder[0].FA.out ),
    .X(net98));
 sky130_fd_sc_hd__buf_1 _431_ (.A(\carry_ripple[2].RA.full_adder[1].FA.out ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _432_ (.A(\carry_ripple[2].RA.full_adder[2].FA.out ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 _433_ (.A(\carry_ripple[2].RA.full_adder[3].FA.out ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 _434_ (.A(\carry_ripple[3].RA.full_adder[0].FA.out ),
    .X(net71));
 sky130_fd_sc_hd__buf_1 _435_ (.A(\carry_ripple[3].RA.full_adder[1].FA.out ),
    .X(net72));
 sky130_fd_sc_hd__buf_1 _436_ (.A(\carry_ripple[3].RA.full_adder[2].FA.out ),
    .X(net73));
 sky130_fd_sc_hd__buf_1 _437_ (.A(\carry_ripple[3].RA.full_adder[3].FA.out ),
    .X(net74));
 sky130_fd_sc_hd__buf_1 _438_ (.A(\carry_ripple[4].RA.full_adder[0].FA.out ),
    .X(net75));
 sky130_fd_sc_hd__buf_1 _439_ (.A(\carry_ripple[4].RA.full_adder[1].FA.out ),
    .X(net76));
 sky130_fd_sc_hd__buf_1 _440_ (.A(\carry_ripple[4].RA.full_adder[2].FA.out ),
    .X(net77));
 sky130_fd_sc_hd__buf_2 _441_ (.A(\carry_ripple[4].RA.full_adder[3].FA.out ),
    .X(net78));
 sky130_fd_sc_hd__buf_1 _442_ (.A(\carry_ripple[5].RA.full_adder[0].FA.out ),
    .X(net80));
 sky130_fd_sc_hd__buf_2 _443_ (.A(\carry_ripple[5].RA.full_adder[1].FA.out ),
    .X(net81));
 sky130_fd_sc_hd__buf_1 _444_ (.A(\carry_ripple[5].RA.full_adder[2].FA.out ),
    .X(net82));
 sky130_fd_sc_hd__buf_1 _445_ (.A(\carry_ripple[5].RA.full_adder[3].FA.out ),
    .X(net83));
 sky130_fd_sc_hd__buf_1 _446_ (.A(\carry_ripple[6].RA.full_adder[0].FA.out ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 _447_ (.A(\carry_ripple[6].RA.full_adder[1].FA.out ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 _448_ (.A(\carry_ripple[6].RA.full_adder[2].FA.out ),
    .X(net86));
 sky130_fd_sc_hd__buf_1 _449_ (.A(\carry_ripple[6].RA.full_adder[3].FA.out ),
    .X(net87));
 sky130_fd_sc_hd__buf_1 _450_ (.A(\carry_ripple[7].RA.full_adder[0].FA.out ),
    .X(net88));
 sky130_fd_sc_hd__buf_1 _451_ (.A(\carry_ripple[7].RA.full_adder[1].FA.out ),
    .X(net89));
 sky130_fd_sc_hd__buf_1 _452_ (.A(\carry_ripple[7].RA.full_adder[2].FA.out ),
    .X(net91));
 sky130_fd_sc_hd__buf_1 _453_ (.A(\carry_ripple[7].RA.full_adder[3].FA.out ),
    .X(net92));
 sky130_fd_sc_hd__buf_2 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(b[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(b[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(b[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(b[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(b[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(b[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(b[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(b[16]),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(b[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(b[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_8 input43 (.A(b[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(b[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(b[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(b[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(b[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(b[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(b[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input50 (.A(b[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(b[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(b[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(b[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(b[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(b[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(b[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(b[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(b[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(b[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(b[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(b[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(b[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(b[8]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(b[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(cin),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_16 output66 (.A(net66),
    .X(cout));
 sky130_fd_sc_hd__clkbuf_16 output67 (.A(net67),
    .X(overflow));
 sky130_fd_sc_hd__clkbuf_16 output68 (.A(net68),
    .X(sum[0]));
 sky130_fd_sc_hd__clkbuf_16 output69 (.A(net69),
    .X(sum[10]));
 sky130_fd_sc_hd__clkbuf_16 output70 (.A(net70),
    .X(sum[11]));
 sky130_fd_sc_hd__clkbuf_16 output71 (.A(net71),
    .X(sum[12]));
 sky130_fd_sc_hd__clkbuf_16 output72 (.A(net72),
    .X(sum[13]));
 sky130_fd_sc_hd__clkbuf_16 output73 (.A(net73),
    .X(sum[14]));
 sky130_fd_sc_hd__clkbuf_16 output74 (.A(net74),
    .X(sum[15]));
 sky130_fd_sc_hd__clkbuf_16 output75 (.A(net75),
    .X(sum[16]));
 sky130_fd_sc_hd__clkbuf_16 output76 (.A(net76),
    .X(sum[17]));
 sky130_fd_sc_hd__clkbuf_16 output77 (.A(net77),
    .X(sum[18]));
 sky130_fd_sc_hd__clkbuf_16 output78 (.A(net78),
    .X(sum[19]));
 sky130_fd_sc_hd__clkbuf_16 output79 (.A(net79),
    .X(sum[1]));
 sky130_fd_sc_hd__clkbuf_16 output80 (.A(net80),
    .X(sum[20]));
 sky130_fd_sc_hd__clkbuf_16 output81 (.A(net81),
    .X(sum[21]));
 sky130_fd_sc_hd__clkbuf_16 output82 (.A(net82),
    .X(sum[22]));
 sky130_fd_sc_hd__clkbuf_16 output83 (.A(net83),
    .X(sum[23]));
 sky130_fd_sc_hd__clkbuf_16 output84 (.A(net84),
    .X(sum[24]));
 sky130_fd_sc_hd__clkbuf_16 output85 (.A(net85),
    .X(sum[25]));
 sky130_fd_sc_hd__clkbuf_16 output86 (.A(net86),
    .X(sum[26]));
 sky130_fd_sc_hd__clkbuf_16 output87 (.A(net87),
    .X(sum[27]));
 sky130_fd_sc_hd__clkbuf_16 output88 (.A(net88),
    .X(sum[28]));
 sky130_fd_sc_hd__clkbuf_16 output89 (.A(net89),
    .X(sum[29]));
 sky130_fd_sc_hd__clkbuf_16 output90 (.A(net90),
    .X(sum[2]));
 sky130_fd_sc_hd__clkbuf_16 output91 (.A(net91),
    .X(sum[30]));
 sky130_fd_sc_hd__clkbuf_16 output92 (.A(net92),
    .X(sum[31]));
 sky130_fd_sc_hd__clkbuf_16 output93 (.A(net93),
    .X(sum[3]));
 sky130_fd_sc_hd__clkbuf_16 output94 (.A(net94),
    .X(sum[4]));
 sky130_fd_sc_hd__clkbuf_16 output95 (.A(net95),
    .X(sum[5]));
 sky130_fd_sc_hd__clkbuf_16 output96 (.A(net96),
    .X(sum[6]));
 sky130_fd_sc_hd__clkbuf_16 output97 (.A(net97),
    .X(sum[7]));
 sky130_fd_sc_hd__clkbuf_16 output98 (.A(net98),
    .X(sum[8]));
 sky130_fd_sc_hd__clkbuf_16 output99 (.A(net99),
    .X(sum[9]));
endmodule
