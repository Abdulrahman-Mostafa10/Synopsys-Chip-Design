module sequential_multiplier_routing(clk,
    reset,
    a,
    b,
    mult);
 input clk;
 input reset;
 input [31:0] a;
 input [31:0] b;
 output [63:0] mult;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \count[4] ;
 wire \count[5] ;
 wire \multiplicand[0] ;
 wire \multiplicand[10] ;
 wire \multiplicand[11] ;
 wire \multiplicand[12] ;
 wire \multiplicand[13] ;
 wire \multiplicand[14] ;
 wire \multiplicand[15] ;
 wire \multiplicand[16] ;
 wire \multiplicand[17] ;
 wire \multiplicand[18] ;
 wire \multiplicand[19] ;
 wire \multiplicand[1] ;
 wire \multiplicand[20] ;
 wire \multiplicand[21] ;
 wire \multiplicand[22] ;
 wire \multiplicand[23] ;
 wire \multiplicand[24] ;
 wire \multiplicand[25] ;
 wire \multiplicand[26] ;
 wire \multiplicand[27] ;
 wire \multiplicand[28] ;
 wire \multiplicand[29] ;
 wire \multiplicand[2] ;
 wire \multiplicand[30] ;
 wire \multiplicand[31] ;
 wire \multiplicand[32] ;
 wire \multiplicand[33] ;
 wire \multiplicand[34] ;
 wire \multiplicand[35] ;
 wire \multiplicand[36] ;
 wire \multiplicand[37] ;
 wire \multiplicand[38] ;
 wire \multiplicand[39] ;
 wire \multiplicand[3] ;
 wire \multiplicand[40] ;
 wire \multiplicand[41] ;
 wire \multiplicand[42] ;
 wire \multiplicand[43] ;
 wire \multiplicand[44] ;
 wire \multiplicand[45] ;
 wire \multiplicand[46] ;
 wire \multiplicand[47] ;
 wire \multiplicand[48] ;
 wire \multiplicand[49] ;
 wire \multiplicand[4] ;
 wire \multiplicand[50] ;
 wire \multiplicand[51] ;
 wire \multiplicand[52] ;
 wire \multiplicand[53] ;
 wire \multiplicand[54] ;
 wire \multiplicand[55] ;
 wire \multiplicand[56] ;
 wire \multiplicand[57] ;
 wire \multiplicand[58] ;
 wire \multiplicand[59] ;
 wire \multiplicand[5] ;
 wire \multiplicand[60] ;
 wire \multiplicand[61] ;
 wire \multiplicand[62] ;
 wire \multiplicand[63] ;
 wire \multiplicand[6] ;
 wire \multiplicand[7] ;
 wire \multiplicand[8] ;
 wire \multiplicand[9] ;
 wire \multiplier[0] ;
 wire \multiplier[10] ;
 wire \multiplier[11] ;
 wire \multiplier[12] ;
 wire \multiplier[13] ;
 wire \multiplier[14] ;
 wire \multiplier[15] ;
 wire \multiplier[16] ;
 wire \multiplier[17] ;
 wire \multiplier[18] ;
 wire \multiplier[19] ;
 wire \multiplier[1] ;
 wire \multiplier[20] ;
 wire \multiplier[21] ;
 wire \multiplier[22] ;
 wire \multiplier[23] ;
 wire \multiplier[24] ;
 wire \multiplier[25] ;
 wire \multiplier[26] ;
 wire \multiplier[27] ;
 wire \multiplier[28] ;
 wire \multiplier[29] ;
 wire \multiplier[2] ;
 wire \multiplier[30] ;
 wire \multiplier[31] ;
 wire \multiplier[3] ;
 wire \multiplier[4] ;
 wire \multiplier[5] ;
 wire \multiplier[6] ;
 wire \multiplier[7] ;
 wire \multiplier[8] ;
 wire \multiplier[9] ;
 wire \product[0] ;
 wire \product[10] ;
 wire \product[11] ;
 wire \product[12] ;
 wire \product[13] ;
 wire \product[14] ;
 wire \product[15] ;
 wire \product[16] ;
 wire \product[17] ;
 wire \product[18] ;
 wire \product[19] ;
 wire \product[1] ;
 wire \product[20] ;
 wire \product[21] ;
 wire \product[22] ;
 wire \product[23] ;
 wire \product[24] ;
 wire \product[25] ;
 wire \product[26] ;
 wire \product[27] ;
 wire \product[28] ;
 wire \product[29] ;
 wire \product[2] ;
 wire \product[30] ;
 wire \product[31] ;
 wire \product[32] ;
 wire \product[33] ;
 wire \product[34] ;
 wire \product[35] ;
 wire \product[36] ;
 wire \product[37] ;
 wire \product[38] ;
 wire \product[39] ;
 wire \product[3] ;
 wire \product[40] ;
 wire \product[41] ;
 wire \product[42] ;
 wire \product[43] ;
 wire \product[44] ;
 wire \product[45] ;
 wire \product[46] ;
 wire \product[47] ;
 wire \product[48] ;
 wire \product[49] ;
 wire \product[4] ;
 wire \product[50] ;
 wire \product[51] ;
 wire \product[52] ;
 wire \product[53] ;
 wire \product[54] ;
 wire \product[55] ;
 wire \product[56] ;
 wire \product[57] ;
 wire \product[58] ;
 wire \product[59] ;
 wire \product[5] ;
 wire \product[60] ;
 wire \product[61] ;
 wire \product[62] ;
 wire \product[63] ;
 wire \product[6] ;
 wire \product[7] ;
 wire \product[8] ;
 wire \product[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_1_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sky130_fd_sc_hd__clkinv_16 _1177_ (.A(net141),
    .Y(_0844_));
 sky130_fd_sc_hd__inv_2 _1178_ (.A(\product[48] ),
    .Y(_0845_));
 sky130_fd_sc_hd__inv_2 _1179_ (.A(\product[46] ),
    .Y(_0846_));
 sky130_fd_sc_hd__inv_2 _1180_ (.A(\product[44] ),
    .Y(_0847_));
 sky130_fd_sc_hd__inv_4 _1181_ (.A(\product[40] ),
    .Y(_0848_));
 sky130_fd_sc_hd__inv_2 _1182_ (.A(\product[34] ),
    .Y(_0849_));
 sky130_fd_sc_hd__inv_4 _1183_ (.A(\product[32] ),
    .Y(_0850_));
 sky130_fd_sc_hd__inv_2 _1184_ (.A(\product[31] ),
    .Y(_0851_));
 sky130_fd_sc_hd__inv_2 _1185_ (.A(\product[28] ),
    .Y(_0852_));
 sky130_fd_sc_hd__inv_2 _1186_ (.A(\product[24] ),
    .Y(_0853_));
 sky130_fd_sc_hd__inv_2 _1187_ (.A(\product[18] ),
    .Y(_0854_));
 sky130_fd_sc_hd__inv_2 _1188_ (.A(\product[16] ),
    .Y(_0855_));
 sky130_fd_sc_hd__clkinv_8 _1189_ (.A(\product[9] ),
    .Y(_0856_));
 sky130_fd_sc_hd__clkinv_8 _1190_ (.A(\product[8] ),
    .Y(_0857_));
 sky130_fd_sc_hd__inv_2 _1191_ (.A(\product[5] ),
    .Y(_0858_));
 sky130_fd_sc_hd__clkinv_16 _1192_ (.A(net65),
    .Y(_0859_));
 sky130_fd_sc_hd__inv_2 _1193_ (.A(net27),
    .Y(_0860_));
 sky130_fd_sc_hd__inv_2 _1194_ (.A(net28),
    .Y(_0861_));
 sky130_fd_sc_hd__inv_2 _1195_ (.A(net29),
    .Y(_0862_));
 sky130_fd_sc_hd__inv_2 _1196_ (.A(net30),
    .Y(_0863_));
 sky130_fd_sc_hd__inv_2 _1197_ (.A(net2),
    .Y(_0864_));
 sky130_fd_sc_hd__inv_2 _1198_ (.A(net5),
    .Y(_0865_));
 sky130_fd_sc_hd__nor2_8 _1199_ (.A(net141),
    .B(net65),
    .Y(_0866_));
 sky130_fd_sc_hd__or2_1 _1200_ (.A(net140),
    .B(net65),
    .X(_0867_));
 sky130_fd_sc_hd__or3_1 _1201_ (.A(net140),
    .B(net65),
    .C(\multiplier[1] ),
    .X(_0868_));
 sky130_fd_sc_hd__nor2_8 _1202_ (.A(net65),
    .B(_0844_),
    .Y(_0869_));
 sky130_fd_sc_hd__nand2_8 _1203_ (.A(_0859_),
    .B(net141),
    .Y(_0870_));
 sky130_fd_sc_hd__o221a_1 _1204_ (.A1(_0859_),
    .A2(net1),
    .B1(_0870_),
    .B2(\multiplier[0] ),
    .C1(_0868_),
    .X(_0000_));
 sky130_fd_sc_hd__a21bo_1 _1205_ (.A1(net25),
    .A2(net1),
    .B1_N(net12),
    .X(_0871_));
 sky130_fd_sc_hd__nand3b_1 _1206_ (.A_N(net12),
    .B(net1),
    .C(net25),
    .Y(_0872_));
 sky130_fd_sc_hd__a21oi_1 _1207_ (.A1(_0871_),
    .A2(_0872_),
    .B1(_0859_),
    .Y(_0873_));
 sky130_fd_sc_hd__a221o_1 _1208_ (.A1(\multiplier[2] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[1] ),
    .C1(_0873_),
    .X(_0001_));
 sky130_fd_sc_hd__o21a_1 _1209_ (.A1(net1),
    .A2(net12),
    .B1(net25),
    .X(_0874_));
 sky130_fd_sc_hd__o21ai_1 _1210_ (.A1(net23),
    .A2(_0874_),
    .B1(net65),
    .Y(_0875_));
 sky130_fd_sc_hd__a21oi_1 _1211_ (.A1(net23),
    .A2(_0874_),
    .B1(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__a221o_1 _1212_ (.A1(\multiplier[3] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[2] ),
    .C1(_0876_),
    .X(_0002_));
 sky130_fd_sc_hd__or3_1 _1213_ (.A(net1),
    .B(net12),
    .C(net23),
    .X(_0877_));
 sky130_fd_sc_hd__o31a_1 _1214_ (.A1(net1),
    .A2(net12),
    .A3(net23),
    .B1(net25),
    .X(_0878_));
 sky130_fd_sc_hd__o21ai_1 _1215_ (.A1(net26),
    .A2(_0878_),
    .B1(net65),
    .Y(_0879_));
 sky130_fd_sc_hd__a21oi_1 _1216_ (.A1(net26),
    .A2(_0878_),
    .B1(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__a221o_1 _1217_ (.A1(\multiplier[4] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[3] ),
    .C1(_0880_),
    .X(_0003_));
 sky130_fd_sc_hd__nor4_1 _1218_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(net26),
    .Y(_0881_));
 sky130_fd_sc_hd__o41a_1 _1219_ (.A1(net1),
    .A2(net12),
    .A3(net23),
    .A4(net26),
    .B1(net25),
    .X(_0882_));
 sky130_fd_sc_hd__a21oi_1 _1220_ (.A1(net27),
    .A2(_0882_),
    .B1(_0859_),
    .Y(_0883_));
 sky130_fd_sc_hd__o21a_1 _1221_ (.A1(net27),
    .A2(_0882_),
    .B1(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__a221o_1 _1222_ (.A1(\multiplier[5] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[4] ),
    .C1(_0884_),
    .X(_0004_));
 sky130_fd_sc_hd__o31a_1 _1223_ (.A1(net26),
    .A2(net27),
    .A3(_0877_),
    .B1(net25),
    .X(_0885_));
 sky130_fd_sc_hd__a21oi_1 _1224_ (.A1(net28),
    .A2(_0885_),
    .B1(_0859_),
    .Y(_0886_));
 sky130_fd_sc_hd__o21a_1 _1225_ (.A1(net28),
    .A2(_0885_),
    .B1(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__a221o_1 _1226_ (.A1(\multiplier[6] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[5] ),
    .C1(_0887_),
    .X(_0005_));
 sky130_fd_sc_hd__o41a_1 _1227_ (.A1(net26),
    .A2(net27),
    .A3(net28),
    .A4(_0877_),
    .B1(net25),
    .X(_0888_));
 sky130_fd_sc_hd__o21ai_1 _1228_ (.A1(net29),
    .A2(_0888_),
    .B1(net65),
    .Y(_0889_));
 sky130_fd_sc_hd__a21oi_1 _1229_ (.A1(net29),
    .A2(_0888_),
    .B1(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__a221o_1 _1230_ (.A1(\multiplier[7] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[6] ),
    .C1(_0890_),
    .X(_0006_));
 sky130_fd_sc_hd__nand4_4 _1231_ (.A(_0881_),
    .B(_0862_),
    .C(_0861_),
    .D(_0860_),
    .Y(_0891_));
 sky130_fd_sc_hd__a21o_1 _1232_ (.A1(_0891_),
    .A2(net25),
    .B1(net30),
    .X(_0892_));
 sky130_fd_sc_hd__nand3_1 _1233_ (.A(_0891_),
    .B(net30),
    .C(net25),
    .Y(_0893_));
 sky130_fd_sc_hd__a22o_1 _1234_ (.A1(\multiplier[8] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[7] ),
    .X(_0894_));
 sky130_fd_sc_hd__a31o_1 _1235_ (.A1(_0892_),
    .A2(_0893_),
    .A3(net65),
    .B1(_0894_),
    .X(_0007_));
 sky130_fd_sc_hd__or2_1 _1236_ (.A(net30),
    .B(_0891_),
    .X(_0895_));
 sky130_fd_sc_hd__o211ai_1 _1237_ (.A1(net30),
    .A2(_0891_),
    .B1(net31),
    .C1(net25),
    .Y(_0896_));
 sky130_fd_sc_hd__a21o_1 _1238_ (.A1(_0895_),
    .A2(net25),
    .B1(net31),
    .X(_0897_));
 sky130_fd_sc_hd__a22o_1 _1239_ (.A1(\multiplier[9] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[8] ),
    .X(_0898_));
 sky130_fd_sc_hd__a31o_1 _1240_ (.A1(_0897_),
    .A2(net65),
    .A3(_0896_),
    .B1(_0898_),
    .X(_0008_));
 sky130_fd_sc_hd__o31a_1 _1241_ (.A1(net30),
    .A2(net31),
    .A3(_0891_),
    .B1(net25),
    .X(_0899_));
 sky130_fd_sc_hd__o21ai_1 _1242_ (.A1(net32),
    .A2(_0899_),
    .B1(net65),
    .Y(_0900_));
 sky130_fd_sc_hd__a21oi_1 _1243_ (.A1(net32),
    .A2(_0899_),
    .B1(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__a221o_1 _1244_ (.A1(\multiplier[10] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[9] ),
    .C1(_0901_),
    .X(_0009_));
 sky130_fd_sc_hd__nor2_1 _1245_ (.A(net31),
    .B(net32),
    .Y(_0902_));
 sky130_fd_sc_hd__o31a_1 _1246_ (.A1(net31),
    .A2(net32),
    .A3(_0895_),
    .B1(net25),
    .X(_0903_));
 sky130_fd_sc_hd__a21oi_1 _1247_ (.A1(net2),
    .A2(_0903_),
    .B1(_0859_),
    .Y(_0904_));
 sky130_fd_sc_hd__o21a_1 _1248_ (.A1(net2),
    .A2(_0903_),
    .B1(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__a221o_1 _1249_ (.A1(\multiplier[11] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[10] ),
    .C1(_0905_),
    .X(_0010_));
 sky130_fd_sc_hd__nand4b_2 _1250_ (.A_N(_0891_),
    .B(_0902_),
    .C(_0863_),
    .D(_0864_),
    .Y(_0906_));
 sky130_fd_sc_hd__o41a_1 _1251_ (.A1(net31),
    .A2(net32),
    .A3(net2),
    .A4(_0895_),
    .B1(net25),
    .X(_0907_));
 sky130_fd_sc_hd__o21ai_1 _1252_ (.A1(net3),
    .A2(_0907_),
    .B1(net65),
    .Y(_0908_));
 sky130_fd_sc_hd__a21oi_1 _1253_ (.A1(net3),
    .A2(_0907_),
    .B1(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__a221o_1 _1254_ (.A1(\multiplier[12] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[11] ),
    .C1(_0909_),
    .X(_0011_));
 sky130_fd_sc_hd__or4b_1 _1255_ (.A(net2),
    .B(net3),
    .C(_0895_),
    .D_N(_0902_),
    .X(_0910_));
 sky130_fd_sc_hd__a21o_1 _1256_ (.A1(_0910_),
    .A2(net25),
    .B1(net4),
    .X(_0911_));
 sky130_fd_sc_hd__o211ai_1 _1257_ (.A1(net3),
    .A2(_0906_),
    .B1(net4),
    .C1(net25),
    .Y(_0912_));
 sky130_fd_sc_hd__a22o_1 _1258_ (.A1(\multiplier[13] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[12] ),
    .X(_0913_));
 sky130_fd_sc_hd__a31o_1 _1259_ (.A1(_0911_),
    .A2(_0912_),
    .A3(net65),
    .B1(_0913_),
    .X(_0012_));
 sky130_fd_sc_hd__nor2_1 _1260_ (.A(net3),
    .B(net4),
    .Y(_0914_));
 sky130_fd_sc_hd__o31a_1 _1261_ (.A1(net3),
    .A2(net4),
    .A3(_0906_),
    .B1(net25),
    .X(_0915_));
 sky130_fd_sc_hd__o21ai_1 _1262_ (.A1(net5),
    .A2(_0915_),
    .B1(net65),
    .Y(_0916_));
 sky130_fd_sc_hd__a21oi_1 _1263_ (.A1(net5),
    .A2(_0915_),
    .B1(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__a221o_1 _1264_ (.A1(\multiplier[14] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[13] ),
    .C1(_0917_),
    .X(_0013_));
 sky130_fd_sc_hd__or4_1 _1265_ (.A(net3),
    .B(net4),
    .C(net5),
    .D(_0906_),
    .X(_0918_));
 sky130_fd_sc_hd__a21oi_1 _1266_ (.A1(_0918_),
    .A2(net25),
    .B1(net6),
    .Y(_0919_));
 sky130_fd_sc_hd__a31o_1 _1267_ (.A1(_0918_),
    .A2(net6),
    .A3(net25),
    .B1(_0859_),
    .X(_0920_));
 sky130_fd_sc_hd__nor2_1 _1268_ (.A(_0919_),
    .B(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__a221o_1 _1269_ (.A1(\multiplier[15] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[14] ),
    .C1(_0921_),
    .X(_0014_));
 sky130_fd_sc_hd__o41a_1 _1270_ (.A1(net4),
    .A2(net5),
    .A3(net6),
    .A4(_0910_),
    .B1(net25),
    .X(_0922_));
 sky130_fd_sc_hd__o21ai_1 _1271_ (.A1(net7),
    .A2(_0922_),
    .B1(net65),
    .Y(_0923_));
 sky130_fd_sc_hd__a21oi_1 _1272_ (.A1(net7),
    .A2(_0922_),
    .B1(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__a221o_1 _1273_ (.A1(\multiplier[16] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[15] ),
    .C1(_0924_),
    .X(_0015_));
 sky130_fd_sc_hd__nor2_1 _1274_ (.A(net6),
    .B(net7),
    .Y(_0925_));
 sky130_fd_sc_hd__nand4b_2 _1275_ (.A_N(_0906_),
    .B(_0914_),
    .C(_0925_),
    .D(_0865_),
    .Y(_0926_));
 sky130_fd_sc_hd__o31a_1 _1276_ (.A1(net6),
    .A2(net7),
    .A3(_0918_),
    .B1(net25),
    .X(_0927_));
 sky130_fd_sc_hd__o21ai_1 _1277_ (.A1(net8),
    .A2(_0927_),
    .B1(net65),
    .Y(_0928_));
 sky130_fd_sc_hd__a21oi_1 _1278_ (.A1(net8),
    .A2(_0927_),
    .B1(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__a221o_1 _1279_ (.A1(\multiplier[17] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[16] ),
    .C1(_0929_),
    .X(_0016_));
 sky130_fd_sc_hd__a211o_1 _1280_ (.A1(net25),
    .A2(net8),
    .B1(net9),
    .C1(_0927_),
    .X(_0930_));
 sky130_fd_sc_hd__o211ai_1 _1281_ (.A1(net8),
    .A2(_0926_),
    .B1(net9),
    .C1(net25),
    .Y(_0931_));
 sky130_fd_sc_hd__a22o_1 _1282_ (.A1(\multiplier[18] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[17] ),
    .X(_0932_));
 sky130_fd_sc_hd__a31o_1 _1283_ (.A1(_0930_),
    .A2(_0931_),
    .A3(net65),
    .B1(_0932_),
    .X(_0017_));
 sky130_fd_sc_hd__nor2_1 _1284_ (.A(net8),
    .B(net9),
    .Y(_0933_));
 sky130_fd_sc_hd__o31a_1 _1285_ (.A1(net8),
    .A2(net9),
    .A3(_0926_),
    .B1(net25),
    .X(_0934_));
 sky130_fd_sc_hd__o21ai_1 _1286_ (.A1(net10),
    .A2(_0934_),
    .B1(net65),
    .Y(_0935_));
 sky130_fd_sc_hd__a21oi_1 _1287_ (.A1(net10),
    .A2(_0934_),
    .B1(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__a221o_1 _1288_ (.A1(\multiplier[19] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[18] ),
    .C1(_0936_),
    .X(_0018_));
 sky130_fd_sc_hd__or4_1 _1289_ (.A(net8),
    .B(net9),
    .C(net10),
    .D(_0926_),
    .X(_0937_));
 sky130_fd_sc_hd__a211o_1 _1290_ (.A1(net25),
    .A2(net10),
    .B1(net11),
    .C1(_0934_),
    .X(_0938_));
 sky130_fd_sc_hd__nand3_1 _1291_ (.A(_0937_),
    .B(net11),
    .C(net25),
    .Y(_0939_));
 sky130_fd_sc_hd__a22o_1 _1292_ (.A1(\multiplier[20] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[19] ),
    .X(_0940_));
 sky130_fd_sc_hd__a31o_1 _1293_ (.A1(_0939_),
    .A2(net65),
    .A3(_0938_),
    .B1(_0940_),
    .X(_0019_));
 sky130_fd_sc_hd__nor2_1 _1294_ (.A(net10),
    .B(net11),
    .Y(_0941_));
 sky130_fd_sc_hd__or4b_1 _1295_ (.A(net10),
    .B(net11),
    .C(_0926_),
    .D_N(_0933_),
    .X(_0942_));
 sky130_fd_sc_hd__and2_1 _1296_ (.A(_0942_),
    .B(net25),
    .X(_0943_));
 sky130_fd_sc_hd__o21ai_1 _1297_ (.A1(net13),
    .A2(_0943_),
    .B1(net65),
    .Y(_0944_));
 sky130_fd_sc_hd__a21oi_1 _1298_ (.A1(net13),
    .A2(_0943_),
    .B1(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__a221o_1 _1299_ (.A1(\multiplier[21] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[20] ),
    .C1(_0945_),
    .X(_0020_));
 sky130_fd_sc_hd__o211ai_1 _1300_ (.A1(net13),
    .A2(_0942_),
    .B1(net14),
    .C1(net25),
    .Y(_0946_));
 sky130_fd_sc_hd__a211o_1 _1301_ (.A1(net25),
    .A2(net13),
    .B1(net14),
    .C1(_0943_),
    .X(_0947_));
 sky130_fd_sc_hd__and3_1 _1302_ (.A(_0947_),
    .B(net65),
    .C(_0946_),
    .X(_0948_));
 sky130_fd_sc_hd__a221o_1 _1303_ (.A1(\multiplier[22] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[21] ),
    .C1(_0948_),
    .X(_0021_));
 sky130_fd_sc_hd__nor2_1 _1304_ (.A(net13),
    .B(net14),
    .Y(_0949_));
 sky130_fd_sc_hd__nand4b_2 _1305_ (.A_N(_0926_),
    .B(_0933_),
    .C(_0941_),
    .D(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__o31a_1 _1306_ (.A1(net13),
    .A2(net14),
    .A3(_0942_),
    .B1(net25),
    .X(_0951_));
 sky130_fd_sc_hd__o21ai_1 _1307_ (.A1(net15),
    .A2(_0951_),
    .B1(net65),
    .Y(_0952_));
 sky130_fd_sc_hd__a21oi_1 _1308_ (.A1(net15),
    .A2(_0951_),
    .B1(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__a221o_1 _1309_ (.A1(\multiplier[23] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[22] ),
    .C1(_0953_),
    .X(_0022_));
 sky130_fd_sc_hd__a211o_1 _1310_ (.A1(net25),
    .A2(net15),
    .B1(net16),
    .C1(_0951_),
    .X(_0954_));
 sky130_fd_sc_hd__o211ai_1 _1311_ (.A1(net15),
    .A2(_0950_),
    .B1(net16),
    .C1(net25),
    .Y(_0955_));
 sky130_fd_sc_hd__a22o_1 _1312_ (.A1(\multiplier[24] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[23] ),
    .X(_0956_));
 sky130_fd_sc_hd__a31o_1 _1313_ (.A1(_0954_),
    .A2(_0955_),
    .A3(net65),
    .B1(_0956_),
    .X(_0023_));
 sky130_fd_sc_hd__or3_1 _1314_ (.A(net15),
    .B(net16),
    .C(_0950_),
    .X(_0957_));
 sky130_fd_sc_hd__o31a_2 _1315_ (.A1(net15),
    .A2(net16),
    .A3(_0950_),
    .B1(net25),
    .X(_0958_));
 sky130_fd_sc_hd__o21ai_1 _1316_ (.A1(net17),
    .A2(_0958_),
    .B1(net65),
    .Y(_0959_));
 sky130_fd_sc_hd__a21oi_1 _1317_ (.A1(net17),
    .A2(_0958_),
    .B1(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__a221o_1 _1318_ (.A1(\multiplier[25] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[24] ),
    .C1(_0960_),
    .X(_0024_));
 sky130_fd_sc_hd__a211o_1 _1319_ (.A1(net25),
    .A2(net17),
    .B1(net18),
    .C1(_0958_),
    .X(_0961_));
 sky130_fd_sc_hd__o211ai_1 _1320_ (.A1(net17),
    .A2(_0957_),
    .B1(net18),
    .C1(net25),
    .Y(_0962_));
 sky130_fd_sc_hd__a22o_1 _1321_ (.A1(\multiplier[26] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[25] ),
    .X(_0963_));
 sky130_fd_sc_hd__a31o_1 _1322_ (.A1(_0962_),
    .A2(net65),
    .A3(_0961_),
    .B1(_0963_),
    .X(_0025_));
 sky130_fd_sc_hd__o21a_1 _1323_ (.A1(net17),
    .A2(net18),
    .B1(net25),
    .X(_0964_));
 sky130_fd_sc_hd__o21ai_1 _1324_ (.A1(_0958_),
    .A2(_0964_),
    .B1(net19),
    .Y(_0965_));
 sky130_fd_sc_hd__or3_1 _1325_ (.A(net19),
    .B(_0958_),
    .C(_0964_),
    .X(_0966_));
 sky130_fd_sc_hd__a22o_1 _1326_ (.A1(\multiplier[27] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[26] ),
    .X(_0967_));
 sky130_fd_sc_hd__a31o_1 _1327_ (.A1(_0966_),
    .A2(net65),
    .A3(_0965_),
    .B1(_0967_),
    .X(_0026_));
 sky130_fd_sc_hd__or3_2 _1328_ (.A(net17),
    .B(net18),
    .C(net19),
    .X(_0968_));
 sky130_fd_sc_hd__a211o_1 _1329_ (.A1(_0968_),
    .A2(net25),
    .B1(net20),
    .C1(_0958_),
    .X(_0969_));
 sky130_fd_sc_hd__o211ai_1 _1330_ (.A1(_0957_),
    .A2(_0968_),
    .B1(net25),
    .C1(net20),
    .Y(_0970_));
 sky130_fd_sc_hd__a22o_1 _1331_ (.A1(\multiplier[28] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[27] ),
    .X(_0971_));
 sky130_fd_sc_hd__a31o_1 _1332_ (.A1(_0970_),
    .A2(net65),
    .A3(_0969_),
    .B1(_0971_),
    .X(_0027_));
 sky130_fd_sc_hd__or4_1 _1333_ (.A(net15),
    .B(net16),
    .C(net20),
    .D(_0968_),
    .X(_0972_));
 sky130_fd_sc_hd__or2_1 _1334_ (.A(_0950_),
    .B(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__nand3_1 _1335_ (.A(_0973_),
    .B(net21),
    .C(net25),
    .Y(_0974_));
 sky130_fd_sc_hd__a21o_1 _1336_ (.A1(_0973_),
    .A2(net25),
    .B1(net21),
    .X(_0975_));
 sky130_fd_sc_hd__a22o_1 _1337_ (.A1(\multiplier[29] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[28] ),
    .X(_0976_));
 sky130_fd_sc_hd__a31o_1 _1338_ (.A1(_0975_),
    .A2(net65),
    .A3(_0974_),
    .B1(_0976_),
    .X(_0028_));
 sky130_fd_sc_hd__or4_1 _1339_ (.A(net20),
    .B(_0968_),
    .C(net21),
    .D(_0957_),
    .X(_0977_));
 sky130_fd_sc_hd__a21o_1 _1340_ (.A1(_0977_),
    .A2(net25),
    .B1(net22),
    .X(_0978_));
 sky130_fd_sc_hd__o211ai_1 _1341_ (.A1(net21),
    .A2(_0973_),
    .B1(net22),
    .C1(net25),
    .Y(_0979_));
 sky130_fd_sc_hd__a22o_1 _1342_ (.A1(\multiplier[30] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[29] ),
    .X(_0980_));
 sky130_fd_sc_hd__a31o_1 _1343_ (.A1(_0978_),
    .A2(_0979_),
    .A3(net65),
    .B1(_0980_),
    .X(_0029_));
 sky130_fd_sc_hd__or3_1 _1344_ (.A(net21),
    .B(net22),
    .C(_0973_),
    .X(_0981_));
 sky130_fd_sc_hd__a21bo_1 _1345_ (.A1(_0981_),
    .A2(net25),
    .B1_N(net24),
    .X(_0982_));
 sky130_fd_sc_hd__nand3b_1 _1346_ (.A_N(net24),
    .B(_0981_),
    .C(net25),
    .Y(_0983_));
 sky130_fd_sc_hd__a21oi_1 _1347_ (.A1(_0982_),
    .A2(_0983_),
    .B1(_0859_),
    .Y(_0984_));
 sky130_fd_sc_hd__a221o_1 _1348_ (.A1(\multiplier[31] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplier[30] ),
    .C1(_0984_),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _1349_ (.A1(net33),
    .A2(net65),
    .B1(\multiplicand[0] ),
    .B2(net136),
    .X(_0031_));
 sky130_fd_sc_hd__or3_1 _1350_ (.A(\count[5] ),
    .B(net65),
    .C(\multiplicand[0] ),
    .X(_0985_));
 sky130_fd_sc_hd__o221a_1 _1351_ (.A1(net142),
    .A2(net44),
    .B1(\multiplicand[1] ),
    .B2(_0870_),
    .C1(_0985_),
    .X(_0032_));
 sky130_fd_sc_hd__or3_1 _1352_ (.A(\count[5] ),
    .B(net65),
    .C(\multiplicand[1] ),
    .X(_0986_));
 sky130_fd_sc_hd__o221a_1 _1353_ (.A1(net142),
    .A2(net55),
    .B1(\multiplicand[2] ),
    .B2(_0870_),
    .C1(_0986_),
    .X(_0033_));
 sky130_fd_sc_hd__or3_1 _1354_ (.A(\count[5] ),
    .B(net65),
    .C(\multiplicand[2] ),
    .X(_0987_));
 sky130_fd_sc_hd__o221a_1 _1355_ (.A1(net142),
    .A2(net58),
    .B1(\multiplicand[3] ),
    .B2(_0870_),
    .C1(_0987_),
    .X(_0034_));
 sky130_fd_sc_hd__or3_1 _1356_ (.A(\count[5] ),
    .B(net65),
    .C(\multiplicand[3] ),
    .X(_0988_));
 sky130_fd_sc_hd__o221a_1 _1357_ (.A1(net142),
    .A2(net59),
    .B1(\multiplicand[4] ),
    .B2(_0870_),
    .C1(_0988_),
    .X(_0035_));
 sky130_fd_sc_hd__or3_1 _1358_ (.A(\count[5] ),
    .B(net65),
    .C(\multiplicand[4] ),
    .X(_0989_));
 sky130_fd_sc_hd__o221a_1 _1359_ (.A1(net142),
    .A2(net60),
    .B1(\multiplicand[5] ),
    .B2(_0870_),
    .C1(_0989_),
    .X(_0036_));
 sky130_fd_sc_hd__or3_1 _1360_ (.A(\count[5] ),
    .B(net65),
    .C(\multiplicand[5] ),
    .X(_0990_));
 sky130_fd_sc_hd__o221a_1 _1361_ (.A1(net142),
    .A2(net61),
    .B1(\multiplicand[6] ),
    .B2(_0870_),
    .C1(_0990_),
    .X(_0037_));
 sky130_fd_sc_hd__or3_1 _1362_ (.A(\count[5] ),
    .B(net65),
    .C(\multiplicand[6] ),
    .X(_0991_));
 sky130_fd_sc_hd__o221a_1 _1363_ (.A1(net142),
    .A2(net62),
    .B1(\multiplicand[7] ),
    .B2(_0870_),
    .C1(_0991_),
    .X(_0038_));
 sky130_fd_sc_hd__or3_1 _1364_ (.A(\count[5] ),
    .B(net65),
    .C(\multiplicand[7] ),
    .X(_0992_));
 sky130_fd_sc_hd__o221a_1 _1365_ (.A1(net142),
    .A2(net63),
    .B1(\multiplicand[8] ),
    .B2(_0870_),
    .C1(_0992_),
    .X(_0039_));
 sky130_fd_sc_hd__or3_1 _1366_ (.A(\count[5] ),
    .B(net65),
    .C(\multiplicand[8] ),
    .X(_0993_));
 sky130_fd_sc_hd__o221a_1 _1367_ (.A1(net142),
    .A2(net64),
    .B1(\multiplicand[9] ),
    .B2(_0870_),
    .C1(_0993_),
    .X(_0040_));
 sky130_fd_sc_hd__or3_1 _1368_ (.A(net139),
    .B(net65),
    .C(\multiplicand[9] ),
    .X(_0994_));
 sky130_fd_sc_hd__o221a_1 _1369_ (.A1(net142),
    .A2(net34),
    .B1(\multiplicand[10] ),
    .B2(_0870_),
    .C1(_0994_),
    .X(_0041_));
 sky130_fd_sc_hd__or3_1 _1370_ (.A(net139),
    .B(net65),
    .C(\multiplicand[10] ),
    .X(_0995_));
 sky130_fd_sc_hd__o221a_1 _1371_ (.A1(net142),
    .A2(net35),
    .B1(\multiplicand[11] ),
    .B2(_0870_),
    .C1(_0995_),
    .X(_0042_));
 sky130_fd_sc_hd__or3_1 _1372_ (.A(net139),
    .B(net65),
    .C(\multiplicand[11] ),
    .X(_0996_));
 sky130_fd_sc_hd__o221a_1 _1373_ (.A1(net142),
    .A2(net36),
    .B1(\multiplicand[12] ),
    .B2(_0870_),
    .C1(_0996_),
    .X(_0043_));
 sky130_fd_sc_hd__or3_1 _1374_ (.A(net139),
    .B(net65),
    .C(\multiplicand[12] ),
    .X(_0997_));
 sky130_fd_sc_hd__o221a_1 _1375_ (.A1(net142),
    .A2(net37),
    .B1(\multiplicand[13] ),
    .B2(_0870_),
    .C1(_0997_),
    .X(_0044_));
 sky130_fd_sc_hd__or3_1 _1376_ (.A(net139),
    .B(net65),
    .C(\multiplicand[13] ),
    .X(_0998_));
 sky130_fd_sc_hd__o221a_1 _1377_ (.A1(net142),
    .A2(net38),
    .B1(\multiplicand[14] ),
    .B2(_0870_),
    .C1(_0998_),
    .X(_0045_));
 sky130_fd_sc_hd__or3_1 _1378_ (.A(net139),
    .B(net65),
    .C(\multiplicand[14] ),
    .X(_0999_));
 sky130_fd_sc_hd__o221a_1 _1379_ (.A1(net142),
    .A2(net39),
    .B1(\multiplicand[15] ),
    .B2(_0870_),
    .C1(_0999_),
    .X(_0046_));
 sky130_fd_sc_hd__or3_1 _1380_ (.A(net139),
    .B(net65),
    .C(\multiplicand[15] ),
    .X(_1000_));
 sky130_fd_sc_hd__o221a_1 _1381_ (.A1(net142),
    .A2(net40),
    .B1(\multiplicand[16] ),
    .B2(_0870_),
    .C1(_1000_),
    .X(_0047_));
 sky130_fd_sc_hd__or3_1 _1382_ (.A(net139),
    .B(net65),
    .C(\multiplicand[16] ),
    .X(_1001_));
 sky130_fd_sc_hd__o221a_1 _1383_ (.A1(net142),
    .A2(net41),
    .B1(\multiplicand[17] ),
    .B2(_0870_),
    .C1(_1001_),
    .X(_0048_));
 sky130_fd_sc_hd__or3_1 _1384_ (.A(net139),
    .B(net65),
    .C(\multiplicand[17] ),
    .X(_1002_));
 sky130_fd_sc_hd__o221a_1 _1385_ (.A1(net142),
    .A2(net42),
    .B1(\multiplicand[18] ),
    .B2(_0870_),
    .C1(_1002_),
    .X(_0049_));
 sky130_fd_sc_hd__or3_1 _1386_ (.A(net139),
    .B(net65),
    .C(\multiplicand[18] ),
    .X(_1003_));
 sky130_fd_sc_hd__o221a_1 _1387_ (.A1(net142),
    .A2(net43),
    .B1(\multiplicand[19] ),
    .B2(_0870_),
    .C1(_1003_),
    .X(_0050_));
 sky130_fd_sc_hd__or3_1 _1388_ (.A(net139),
    .B(net65),
    .C(\multiplicand[19] ),
    .X(_1004_));
 sky130_fd_sc_hd__o221a_1 _1389_ (.A1(net142),
    .A2(net45),
    .B1(\multiplicand[20] ),
    .B2(_0870_),
    .C1(_1004_),
    .X(_0051_));
 sky130_fd_sc_hd__or3_1 _1390_ (.A(net139),
    .B(net65),
    .C(\multiplicand[20] ),
    .X(_1005_));
 sky130_fd_sc_hd__o221a_1 _1391_ (.A1(net142),
    .A2(net46),
    .B1(\multiplicand[21] ),
    .B2(_0870_),
    .C1(_1005_),
    .X(_0052_));
 sky130_fd_sc_hd__or3_1 _1392_ (.A(net139),
    .B(net65),
    .C(\multiplicand[21] ),
    .X(_1006_));
 sky130_fd_sc_hd__o221a_1 _1393_ (.A1(net142),
    .A2(net47),
    .B1(\multiplicand[22] ),
    .B2(_0870_),
    .C1(_1006_),
    .X(_0053_));
 sky130_fd_sc_hd__or3_1 _1394_ (.A(net139),
    .B(net65),
    .C(\multiplicand[22] ),
    .X(_1007_));
 sky130_fd_sc_hd__o221a_1 _1395_ (.A1(net142),
    .A2(net48),
    .B1(\multiplicand[23] ),
    .B2(_0870_),
    .C1(_1007_),
    .X(_0054_));
 sky130_fd_sc_hd__or3_1 _1396_ (.A(net139),
    .B(net65),
    .C(\multiplicand[23] ),
    .X(_1008_));
 sky130_fd_sc_hd__o221a_1 _1397_ (.A1(net142),
    .A2(net49),
    .B1(\multiplicand[24] ),
    .B2(_0870_),
    .C1(_1008_),
    .X(_0055_));
 sky130_fd_sc_hd__or3_1 _1398_ (.A(net139),
    .B(net65),
    .C(\multiplicand[24] ),
    .X(_1009_));
 sky130_fd_sc_hd__o221a_1 _1399_ (.A1(net142),
    .A2(net50),
    .B1(\multiplicand[25] ),
    .B2(_0870_),
    .C1(_1009_),
    .X(_0056_));
 sky130_fd_sc_hd__or3_1 _1400_ (.A(net139),
    .B(net65),
    .C(\multiplicand[25] ),
    .X(_1010_));
 sky130_fd_sc_hd__o221a_1 _1401_ (.A1(net142),
    .A2(net51),
    .B1(\multiplicand[26] ),
    .B2(_0870_),
    .C1(_1010_),
    .X(_0057_));
 sky130_fd_sc_hd__or3_1 _1402_ (.A(net139),
    .B(net65),
    .C(\multiplicand[26] ),
    .X(_1011_));
 sky130_fd_sc_hd__o221a_1 _1403_ (.A1(net142),
    .A2(net52),
    .B1(\multiplicand[27] ),
    .B2(_0870_),
    .C1(_1011_),
    .X(_0058_));
 sky130_fd_sc_hd__or3_1 _1404_ (.A(net139),
    .B(net65),
    .C(\multiplicand[27] ),
    .X(_1012_));
 sky130_fd_sc_hd__o221a_1 _1405_ (.A1(net142),
    .A2(net53),
    .B1(\multiplicand[28] ),
    .B2(_0870_),
    .C1(_1012_),
    .X(_0059_));
 sky130_fd_sc_hd__or3_1 _1406_ (.A(net139),
    .B(net65),
    .C(\multiplicand[28] ),
    .X(_1013_));
 sky130_fd_sc_hd__o221a_1 _1407_ (.A1(net142),
    .A2(net54),
    .B1(\multiplicand[29] ),
    .B2(_0870_),
    .C1(_1013_),
    .X(_0060_));
 sky130_fd_sc_hd__or3_1 _1408_ (.A(net139),
    .B(net65),
    .C(\multiplicand[29] ),
    .X(_1014_));
 sky130_fd_sc_hd__o221a_1 _1409_ (.A1(net142),
    .A2(net56),
    .B1(\multiplicand[30] ),
    .B2(_0870_),
    .C1(_1014_),
    .X(_0061_));
 sky130_fd_sc_hd__and2_4 _1410_ (.A(net65),
    .B(net57),
    .X(_1015_));
 sky130_fd_sc_hd__a221o_1 _1411_ (.A1(\multiplicand[30] ),
    .A2(net138),
    .B1(net136),
    .B2(\multiplicand[31] ),
    .C1(_1015_),
    .X(_0062_));
 sky130_fd_sc_hd__a221o_1 _1412_ (.A1(\multiplicand[31] ),
    .A2(net138),
    .B1(net136),
    .B2(\multiplicand[32] ),
    .C1(_1015_),
    .X(_0063_));
 sky130_fd_sc_hd__a221o_1 _1413_ (.A1(\multiplicand[32] ),
    .A2(_0866_),
    .B1(net136),
    .B2(\multiplicand[33] ),
    .C1(_1015_),
    .X(_0064_));
 sky130_fd_sc_hd__a221o_1 _1414_ (.A1(\multiplicand[33] ),
    .A2(_0866_),
    .B1(net136),
    .B2(\multiplicand[34] ),
    .C1(_1015_),
    .X(_0065_));
 sky130_fd_sc_hd__a221o_1 _1415_ (.A1(\multiplicand[34] ),
    .A2(_0866_),
    .B1(net136),
    .B2(\multiplicand[35] ),
    .C1(_1015_),
    .X(_0066_));
 sky130_fd_sc_hd__a221o_1 _1416_ (.A1(\multiplicand[35] ),
    .A2(_0866_),
    .B1(net136),
    .B2(\multiplicand[36] ),
    .C1(_1015_),
    .X(_0067_));
 sky130_fd_sc_hd__a221o_1 _1417_ (.A1(\multiplicand[36] ),
    .A2(_0866_),
    .B1(net136),
    .B2(\multiplicand[37] ),
    .C1(_1015_),
    .X(_0068_));
 sky130_fd_sc_hd__a221o_1 _1418_ (.A1(\multiplicand[37] ),
    .A2(_0866_),
    .B1(net136),
    .B2(\multiplicand[38] ),
    .C1(_1015_),
    .X(_0069_));
 sky130_fd_sc_hd__a221o_1 _1419_ (.A1(\multiplicand[38] ),
    .A2(_0866_),
    .B1(net136),
    .B2(\multiplicand[39] ),
    .C1(_1015_),
    .X(_0070_));
 sky130_fd_sc_hd__a221o_1 _1420_ (.A1(\multiplicand[39] ),
    .A2(_0866_),
    .B1(net136),
    .B2(\multiplicand[40] ),
    .C1(_1015_),
    .X(_0071_));
 sky130_fd_sc_hd__a221o_1 _1421_ (.A1(\multiplicand[40] ),
    .A2(_0866_),
    .B1(net136),
    .B2(\multiplicand[41] ),
    .C1(_1015_),
    .X(_0072_));
 sky130_fd_sc_hd__a221o_1 _1422_ (.A1(\multiplicand[41] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[42] ),
    .C1(_1015_),
    .X(_0073_));
 sky130_fd_sc_hd__a221o_1 _1423_ (.A1(\multiplicand[42] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[43] ),
    .C1(_1015_),
    .X(_0074_));
 sky130_fd_sc_hd__a221o_1 _1424_ (.A1(\multiplicand[43] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[44] ),
    .C1(_1015_),
    .X(_0075_));
 sky130_fd_sc_hd__a221o_1 _1425_ (.A1(\multiplicand[44] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[45] ),
    .C1(_1015_),
    .X(_0076_));
 sky130_fd_sc_hd__a221o_1 _1426_ (.A1(\multiplicand[45] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[46] ),
    .C1(_1015_),
    .X(_0077_));
 sky130_fd_sc_hd__a221o_1 _1427_ (.A1(\multiplicand[46] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[47] ),
    .C1(_1015_),
    .X(_0078_));
 sky130_fd_sc_hd__a221o_1 _1428_ (.A1(\multiplicand[47] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[48] ),
    .C1(_1015_),
    .X(_0079_));
 sky130_fd_sc_hd__a221o_1 _1429_ (.A1(\multiplicand[48] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[49] ),
    .C1(_1015_),
    .X(_0080_));
 sky130_fd_sc_hd__a221o_1 _1430_ (.A1(\multiplicand[49] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[50] ),
    .C1(_1015_),
    .X(_0081_));
 sky130_fd_sc_hd__a221o_1 _1431_ (.A1(\multiplicand[50] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[51] ),
    .C1(_1015_),
    .X(_0082_));
 sky130_fd_sc_hd__a221o_1 _1432_ (.A1(\multiplicand[51] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[52] ),
    .C1(_1015_),
    .X(_0083_));
 sky130_fd_sc_hd__a221o_1 _1433_ (.A1(\multiplicand[52] ),
    .A2(_0866_),
    .B1(_0869_),
    .B2(\multiplicand[53] ),
    .C1(_1015_),
    .X(_0084_));
 sky130_fd_sc_hd__a221o_1 _1434_ (.A1(\multiplicand[53] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplicand[54] ),
    .C1(_1015_),
    .X(_0085_));
 sky130_fd_sc_hd__a221o_1 _1435_ (.A1(\multiplicand[54] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplicand[55] ),
    .C1(_1015_),
    .X(_0086_));
 sky130_fd_sc_hd__a221o_1 _1436_ (.A1(\multiplicand[55] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplicand[56] ),
    .C1(_1015_),
    .X(_0087_));
 sky130_fd_sc_hd__a221o_1 _1437_ (.A1(\multiplicand[56] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplicand[57] ),
    .C1(_1015_),
    .X(_0088_));
 sky130_fd_sc_hd__a221o_1 _1438_ (.A1(\multiplicand[57] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplicand[58] ),
    .C1(_1015_),
    .X(_0089_));
 sky130_fd_sc_hd__a221o_1 _1439_ (.A1(\multiplicand[58] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplicand[59] ),
    .C1(_1015_),
    .X(_0090_));
 sky130_fd_sc_hd__a221o_1 _1440_ (.A1(\multiplicand[59] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplicand[60] ),
    .C1(_1015_),
    .X(_0091_));
 sky130_fd_sc_hd__a221o_1 _1441_ (.A1(\multiplicand[60] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplicand[61] ),
    .C1(_1015_),
    .X(_0092_));
 sky130_fd_sc_hd__a221o_1 _1442_ (.A1(\multiplicand[61] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplicand[62] ),
    .C1(_1015_),
    .X(_0093_));
 sky130_fd_sc_hd__a221o_1 _1443_ (.A1(\multiplicand[62] ),
    .A2(net137),
    .B1(net135),
    .B2(\multiplicand[63] ),
    .C1(_1015_),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _1444_ (.A1(net66),
    .A2(net138),
    .B1(net136),
    .B2(\product[0] ),
    .X(_0095_));
 sky130_fd_sc_hd__nand2_1 _1445_ (.A(\product[0] ),
    .B(net25),
    .Y(_1016_));
 sky130_fd_sc_hd__nor2_1 _1446_ (.A(\product[1] ),
    .B(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__a21o_1 _1447_ (.A1(_1016_),
    .A2(\product[1] ),
    .B1(_0844_),
    .X(_1018_));
 sky130_fd_sc_hd__o221a_1 _1448_ (.A1(\count[5] ),
    .A2(net77),
    .B1(_1017_),
    .B2(_1018_),
    .C1(net142),
    .X(_0096_));
 sky130_fd_sc_hd__or2_1 _1449_ (.A(\product[1] ),
    .B(\product[0] ),
    .X(_1019_));
 sky130_fd_sc_hd__o21ai_1 _1450_ (.A1(\product[1] ),
    .A2(\product[0] ),
    .B1(net25),
    .Y(_1020_));
 sky130_fd_sc_hd__a21oi_1 _1451_ (.A1(_1020_),
    .A2(\product[2] ),
    .B1(_0844_),
    .Y(_1021_));
 sky130_fd_sc_hd__o21ai_1 _1452_ (.A1(\product[2] ),
    .A2(_1020_),
    .B1(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__o211a_1 _1453_ (.A1(\count[5] ),
    .A2(net88),
    .B1(net142),
    .C1(_1022_),
    .X(_0097_));
 sky130_fd_sc_hd__nor3_2 _1454_ (.A(\product[2] ),
    .B(\product[1] ),
    .C(\product[0] ),
    .Y(_1023_));
 sky130_fd_sc_hd__or3_1 _1455_ (.A(\product[2] ),
    .B(\product[1] ),
    .C(\product[0] ),
    .X(_1024_));
 sky130_fd_sc_hd__o21ai_1 _1456_ (.A1(\product[2] ),
    .A2(_1019_),
    .B1(net25),
    .Y(_1025_));
 sky130_fd_sc_hd__a21oi_1 _1457_ (.A1(_1025_),
    .A2(\product[3] ),
    .B1(_0844_),
    .Y(_1026_));
 sky130_fd_sc_hd__o21ai_1 _1458_ (.A1(\product[3] ),
    .A2(_1025_),
    .B1(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__o211a_1 _1459_ (.A1(\count[5] ),
    .A2(net99),
    .B1(net142),
    .C1(_1027_),
    .X(_0098_));
 sky130_fd_sc_hd__o21ai_1 _1460_ (.A1(\product[3] ),
    .A2(_1024_),
    .B1(net25),
    .Y(_1028_));
 sky130_fd_sc_hd__a21oi_1 _1461_ (.A1(_1028_),
    .A2(\product[4] ),
    .B1(_0844_),
    .Y(_1029_));
 sky130_fd_sc_hd__o21ai_1 _1462_ (.A1(\product[4] ),
    .A2(_1028_),
    .B1(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__o211a_1 _1463_ (.A1(\count[5] ),
    .A2(net110),
    .B1(net142),
    .C1(_1030_),
    .X(_0099_));
 sky130_fd_sc_hd__nor2_1 _1464_ (.A(\product[4] ),
    .B(\product[3] ),
    .Y(_1031_));
 sky130_fd_sc_hd__or4_1 _1465_ (.A(\product[4] ),
    .B(\product[3] ),
    .C(\product[2] ),
    .D(_1019_),
    .X(_1032_));
 sky130_fd_sc_hd__a21oi_1 _1466_ (.A1(_1032_),
    .A2(net25),
    .B1(_0858_),
    .Y(_1033_));
 sky130_fd_sc_hd__a31o_1 _1467_ (.A1(_0858_),
    .A2(_1032_),
    .A3(net25),
    .B1(_0844_),
    .X(_1034_));
 sky130_fd_sc_hd__o221a_1 _1468_ (.A1(\count[5] ),
    .A2(net121),
    .B1(_1033_),
    .B2(_1034_),
    .C1(net142),
    .X(_0100_));
 sky130_fd_sc_hd__or4_1 _1469_ (.A(\product[5] ),
    .B(\product[4] ),
    .C(\product[3] ),
    .D(_1024_),
    .X(_1035_));
 sky130_fd_sc_hd__o21ai_1 _1470_ (.A1(\product[5] ),
    .A2(_1032_),
    .B1(net25),
    .Y(_1036_));
 sky130_fd_sc_hd__a21oi_1 _1471_ (.A1(_1036_),
    .A2(\product[6] ),
    .B1(_0844_),
    .Y(_1037_));
 sky130_fd_sc_hd__o21ai_1 _1472_ (.A1(\product[6] ),
    .A2(_1036_),
    .B1(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__o211a_1 _1473_ (.A1(\count[5] ),
    .A2(net126),
    .B1(net142),
    .C1(_1038_),
    .X(_0101_));
 sky130_fd_sc_hd__nor2_1 _1474_ (.A(\product[6] ),
    .B(\product[5] ),
    .Y(_1039_));
 sky130_fd_sc_hd__o21ai_1 _1475_ (.A1(\product[6] ),
    .A2(_1035_),
    .B1(net25),
    .Y(_1040_));
 sky130_fd_sc_hd__nor2_1 _1476_ (.A(\product[7] ),
    .B(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__a21o_1 _1477_ (.A1(_1040_),
    .A2(\product[7] ),
    .B1(_0844_),
    .X(_1042_));
 sky130_fd_sc_hd__o221a_1 _1478_ (.A1(\count[5] ),
    .A2(net127),
    .B1(_1041_),
    .B2(_1042_),
    .C1(net142),
    .X(_0102_));
 sky130_fd_sc_hd__nand4b_4 _1479_ (.A_N(\product[7] ),
    .B(_1023_),
    .C(_1031_),
    .D(_1039_),
    .Y(_1043_));
 sky130_fd_sc_hd__a21oi_1 _1480_ (.A1(_1043_),
    .A2(net25),
    .B1(_0857_),
    .Y(_1044_));
 sky130_fd_sc_hd__a31o_1 _1481_ (.A1(_0857_),
    .A2(_1043_),
    .A3(net25),
    .B1(_0844_),
    .X(_1045_));
 sky130_fd_sc_hd__o221a_1 _1482_ (.A1(\count[5] ),
    .A2(net128),
    .B1(_1044_),
    .B2(_1045_),
    .C1(net142),
    .X(_0103_));
 sky130_fd_sc_hd__o41a_1 _1483_ (.A1(\product[8] ),
    .A2(\product[7] ),
    .A3(\product[6] ),
    .A4(_1035_),
    .B1(net25),
    .X(_1046_));
 sky130_fd_sc_hd__o211a_1 _1484_ (.A1(\product[8] ),
    .A2(_1043_),
    .B1(net25),
    .C1(_0856_),
    .X(_1047_));
 sky130_fd_sc_hd__o21ai_1 _1485_ (.A1(_0856_),
    .A2(_1046_),
    .B1(\count[5] ),
    .Y(_1048_));
 sky130_fd_sc_hd__o221a_1 _1486_ (.A1(\count[5] ),
    .A2(net129),
    .B1(_1047_),
    .B2(_1048_),
    .C1(net142),
    .X(_0104_));
 sky130_fd_sc_hd__or3_4 _1487_ (.A(\product[9] ),
    .B(\product[8] ),
    .C(_1043_),
    .X(_1049_));
 sky130_fd_sc_hd__a21oi_1 _1488_ (.A1(_1049_),
    .A2(net25),
    .B1(\product[10] ),
    .Y(_1050_));
 sky130_fd_sc_hd__a31o_1 _1489_ (.A1(_1049_),
    .A2(net25),
    .A3(\product[10] ),
    .B1(_0870_),
    .X(_1051_));
 sky130_fd_sc_hd__a2bb2o_1 _1490_ (.A1_N(_1050_),
    .A2_N(_1051_),
    .B1(net67),
    .B2(net138),
    .X(_0105_));
 sky130_fd_sc_hd__o21ai_1 _1491_ (.A1(\product[10] ),
    .A2(_1049_),
    .B1(net25),
    .Y(_1052_));
 sky130_fd_sc_hd__a21oi_1 _1492_ (.A1(\product[11] ),
    .A2(_1052_),
    .B1(_0844_),
    .Y(_1053_));
 sky130_fd_sc_hd__o21ai_2 _1493_ (.A1(\product[11] ),
    .A2(_1052_),
    .B1(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__o211a_1 _1494_ (.A1(net139),
    .A2(net68),
    .B1(net142),
    .C1(_1054_),
    .X(_0106_));
 sky130_fd_sc_hd__nor2_1 _1495_ (.A(\product[11] ),
    .B(\product[10] ),
    .Y(_1055_));
 sky130_fd_sc_hd__nor4b_4 _1496_ (.A(\product[9] ),
    .B(\product[8] ),
    .C(_1043_),
    .D_N(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__o31ai_2 _1497_ (.A1(\product[11] ),
    .A2(\product[10] ),
    .A3(_1049_),
    .B1(net25),
    .Y(_1057_));
 sky130_fd_sc_hd__o21ai_1 _1498_ (.A1(\product[12] ),
    .A2(_1057_),
    .B1(net139),
    .Y(_1058_));
 sky130_fd_sc_hd__a21o_1 _1499_ (.A1(\product[12] ),
    .A2(_1057_),
    .B1(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__o211a_1 _1500_ (.A1(net139),
    .A2(net69),
    .B1(net142),
    .C1(_1059_),
    .X(_0107_));
 sky130_fd_sc_hd__o41a_1 _1501_ (.A1(\product[12] ),
    .A2(\product[11] ),
    .A3(\product[10] ),
    .A4(_1049_),
    .B1(net25),
    .X(_1060_));
 sky130_fd_sc_hd__o21ai_1 _1502_ (.A1(\product[13] ),
    .A2(_1060_),
    .B1(net136),
    .Y(_1061_));
 sky130_fd_sc_hd__a21oi_2 _1503_ (.A1(\product[13] ),
    .A2(_1060_),
    .B1(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__a31o_1 _1504_ (.A1(_0844_),
    .A2(net70),
    .A3(net142),
    .B1(_1062_),
    .X(_0108_));
 sky130_fd_sc_hd__nor2_2 _1505_ (.A(\product[13] ),
    .B(\product[12] ),
    .Y(_1063_));
 sky130_fd_sc_hd__or4b_2 _1506_ (.A(\product[13] ),
    .B(\product[12] ),
    .C(_1049_),
    .D_N(_1055_),
    .X(_1064_));
 sky130_fd_sc_hd__nand2_1 _1507_ (.A(_1064_),
    .B(net25),
    .Y(_1065_));
 sky130_fd_sc_hd__a21oi_1 _1508_ (.A1(_1065_),
    .A2(\product[14] ),
    .B1(_0844_),
    .Y(_1066_));
 sky130_fd_sc_hd__o21ai_1 _1509_ (.A1(\product[14] ),
    .A2(_1065_),
    .B1(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__o211a_1 _1510_ (.A1(net139),
    .A2(net71),
    .B1(net142),
    .C1(_1067_),
    .X(_0109_));
 sky130_fd_sc_hd__o21ai_1 _1511_ (.A1(\product[14] ),
    .A2(_1064_),
    .B1(net25),
    .Y(_1068_));
 sky130_fd_sc_hd__o21ai_1 _1512_ (.A1(\product[15] ),
    .A2(_1068_),
    .B1(net139),
    .Y(_1069_));
 sky130_fd_sc_hd__a21o_1 _1513_ (.A1(\product[15] ),
    .A2(_1068_),
    .B1(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__o211a_1 _1514_ (.A1(net139),
    .A2(net72),
    .B1(net142),
    .C1(_1070_),
    .X(_0110_));
 sky130_fd_sc_hd__nor2_2 _1515_ (.A(\product[15] ),
    .B(\product[14] ),
    .Y(_1071_));
 sky130_fd_sc_hd__nand3_4 _1516_ (.A(_1056_),
    .B(_1063_),
    .C(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__a21oi_1 _1517_ (.A1(_1072_),
    .A2(net25),
    .B1(_0855_),
    .Y(_1073_));
 sky130_fd_sc_hd__a31o_1 _1518_ (.A1(_0855_),
    .A2(_1072_),
    .A3(net25),
    .B1(_0844_),
    .X(_1074_));
 sky130_fd_sc_hd__o221a_1 _1519_ (.A1(net139),
    .A2(net73),
    .B1(_1073_),
    .B2(_1074_),
    .C1(net142),
    .X(_0111_));
 sky130_fd_sc_hd__o21ai_1 _1520_ (.A1(\product[16] ),
    .A2(_1072_),
    .B1(net25),
    .Y(_1075_));
 sky130_fd_sc_hd__o21ai_1 _1521_ (.A1(\product[17] ),
    .A2(_1075_),
    .B1(net139),
    .Y(_1076_));
 sky130_fd_sc_hd__a21o_1 _1522_ (.A1(\product[17] ),
    .A2(_1075_),
    .B1(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__o211a_1 _1523_ (.A1(net139),
    .A2(net74),
    .B1(net142),
    .C1(_1077_),
    .X(_0112_));
 sky130_fd_sc_hd__or3_2 _1524_ (.A(\product[17] ),
    .B(\product[16] ),
    .C(_1072_),
    .X(_1078_));
 sky130_fd_sc_hd__a21oi_1 _1525_ (.A1(_1078_),
    .A2(net25),
    .B1(_0854_),
    .Y(_1079_));
 sky130_fd_sc_hd__a31o_1 _1526_ (.A1(_0854_),
    .A2(_1078_),
    .A3(net25),
    .B1(_0844_),
    .X(_1080_));
 sky130_fd_sc_hd__o221a_1 _1527_ (.A1(net139),
    .A2(net75),
    .B1(_1079_),
    .B2(_1080_),
    .C1(net142),
    .X(_0113_));
 sky130_fd_sc_hd__o21ai_1 _1528_ (.A1(\product[18] ),
    .A2(_1078_),
    .B1(net25),
    .Y(_1081_));
 sky130_fd_sc_hd__o21ai_1 _1529_ (.A1(\product[19] ),
    .A2(_1081_),
    .B1(net139),
    .Y(_1082_));
 sky130_fd_sc_hd__a21o_1 _1530_ (.A1(\product[19] ),
    .A2(_1081_),
    .B1(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__o211a_1 _1531_ (.A1(net139),
    .A2(net76),
    .B1(net142),
    .C1(_1083_),
    .X(_0114_));
 sky130_fd_sc_hd__or3_1 _1532_ (.A(\product[19] ),
    .B(\product[18] ),
    .C(_1078_),
    .X(_1084_));
 sky130_fd_sc_hd__nand2_1 _1533_ (.A(_1084_),
    .B(net25),
    .Y(_1085_));
 sky130_fd_sc_hd__o21ai_1 _1534_ (.A1(\product[20] ),
    .A2(_1085_),
    .B1(net139),
    .Y(_1086_));
 sky130_fd_sc_hd__a21o_1 _1535_ (.A1(\product[20] ),
    .A2(_1085_),
    .B1(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__o211a_1 _1536_ (.A1(net139),
    .A2(net78),
    .B1(net142),
    .C1(_1087_),
    .X(_0115_));
 sky130_fd_sc_hd__o21ai_1 _1537_ (.A1(\product[20] ),
    .A2(_1084_),
    .B1(net25),
    .Y(_1088_));
 sky130_fd_sc_hd__o21ai_1 _1538_ (.A1(\product[21] ),
    .A2(_1088_),
    .B1(net139),
    .Y(_1089_));
 sky130_fd_sc_hd__a21o_1 _1539_ (.A1(\product[21] ),
    .A2(_1088_),
    .B1(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__o211a_1 _1540_ (.A1(net139),
    .A2(net79),
    .B1(net142),
    .C1(_1090_),
    .X(_0116_));
 sky130_fd_sc_hd__or3_2 _1541_ (.A(\product[20] ),
    .B(\product[19] ),
    .C(\product[18] ),
    .X(_1091_));
 sky130_fd_sc_hd__o31ai_1 _1542_ (.A1(_1091_),
    .A2(\product[21] ),
    .A3(_1078_),
    .B1(net25),
    .Y(_1092_));
 sky130_fd_sc_hd__o21ai_1 _1543_ (.A1(\product[22] ),
    .A2(_1092_),
    .B1(net139),
    .Y(_1093_));
 sky130_fd_sc_hd__a21o_1 _1544_ (.A1(\product[22] ),
    .A2(_1092_),
    .B1(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__o211a_1 _1545_ (.A1(net139),
    .A2(net80),
    .B1(net142),
    .C1(_1094_),
    .X(_0117_));
 sky130_fd_sc_hd__or4_1 _1546_ (.A(\product[22] ),
    .B(\product[21] ),
    .C(\product[20] ),
    .D(_1084_),
    .X(_1095_));
 sky130_fd_sc_hd__nand3b_1 _1547_ (.A_N(\product[23] ),
    .B(_1095_),
    .C(net25),
    .Y(_1096_));
 sky130_fd_sc_hd__a21bo_1 _1548_ (.A1(_1095_),
    .A2(net25),
    .B1_N(\product[23] ),
    .X(_1097_));
 sky130_fd_sc_hd__nor2_1 _1549_ (.A(net139),
    .B(net81),
    .Y(_1098_));
 sky130_fd_sc_hd__a311oi_1 _1550_ (.A1(_1097_),
    .A2(net139),
    .A3(_1096_),
    .B1(_1098_),
    .C1(net65),
    .Y(_0118_));
 sky130_fd_sc_hd__or4_1 _1551_ (.A(\product[23] ),
    .B(\product[22] ),
    .C(\product[17] ),
    .D(\product[16] ),
    .X(_1099_));
 sky130_fd_sc_hd__nor3_4 _1552_ (.A(\product[21] ),
    .B(_1091_),
    .C(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__nand4_4 _1553_ (.A(_1056_),
    .B(_1063_),
    .C(_1071_),
    .D(_1100_),
    .Y(_1101_));
 sky130_fd_sc_hd__a21oi_1 _1554_ (.A1(_1101_),
    .A2(net25),
    .B1(_0853_),
    .Y(_1102_));
 sky130_fd_sc_hd__a31o_1 _1555_ (.A1(_0853_),
    .A2(_1101_),
    .A3(net25),
    .B1(_0844_),
    .X(_1103_));
 sky130_fd_sc_hd__o221a_1 _1556_ (.A1(net139),
    .A2(net82),
    .B1(_1102_),
    .B2(_1103_),
    .C1(net142),
    .X(_0119_));
 sky130_fd_sc_hd__o21ai_1 _1557_ (.A1(\product[24] ),
    .A2(_1101_),
    .B1(net25),
    .Y(_1104_));
 sky130_fd_sc_hd__o21ai_1 _1558_ (.A1(\product[25] ),
    .A2(_1104_),
    .B1(net139),
    .Y(_1105_));
 sky130_fd_sc_hd__a21o_4 _1559_ (.A1(\product[25] ),
    .A2(_1104_),
    .B1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__o211a_1 _1560_ (.A1(net141),
    .A2(net83),
    .B1(_0859_),
    .C1(_1106_),
    .X(_0120_));
 sky130_fd_sc_hd__o31ai_1 _1561_ (.A1(\product[25] ),
    .A2(\product[24] ),
    .A3(_1101_),
    .B1(net25),
    .Y(_1107_));
 sky130_fd_sc_hd__o21ai_1 _1562_ (.A1(\product[26] ),
    .A2(_1107_),
    .B1(net139),
    .Y(_1108_));
 sky130_fd_sc_hd__a21o_1 _1563_ (.A1(\product[26] ),
    .A2(_1107_),
    .B1(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__o211a_1 _1564_ (.A1(net139),
    .A2(net84),
    .B1(net142),
    .C1(_1109_),
    .X(_0121_));
 sky130_fd_sc_hd__o41ai_2 _1565_ (.A1(\product[26] ),
    .A2(\product[25] ),
    .A3(\product[24] ),
    .A4(_1101_),
    .B1(net25),
    .Y(_1110_));
 sky130_fd_sc_hd__o21ai_1 _1566_ (.A1(\product[27] ),
    .A2(_1110_),
    .B1(net139),
    .Y(_1111_));
 sky130_fd_sc_hd__a21o_4 _1567_ (.A1(\product[27] ),
    .A2(_1110_),
    .B1(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__o211a_1 _1568_ (.A1(net141),
    .A2(net85),
    .B1(_0859_),
    .C1(_1112_),
    .X(_0122_));
 sky130_fd_sc_hd__nor4_4 _1569_ (.A(\product[27] ),
    .B(\product[26] ),
    .C(\product[25] ),
    .D(\product[24] ),
    .Y(_1113_));
 sky130_fd_sc_hd__nand3b_2 _1570_ (.A_N(_1072_),
    .B(_1100_),
    .C(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__a21oi_1 _1571_ (.A1(_1114_),
    .A2(net25),
    .B1(_0852_),
    .Y(_1115_));
 sky130_fd_sc_hd__a31o_1 _1572_ (.A1(_0852_),
    .A2(_1114_),
    .A3(net25),
    .B1(_0844_),
    .X(_1116_));
 sky130_fd_sc_hd__o221a_1 _1573_ (.A1(net139),
    .A2(net86),
    .B1(_1115_),
    .B2(_1116_),
    .C1(net142),
    .X(_0123_));
 sky130_fd_sc_hd__o21a_1 _1574_ (.A1(\product[28] ),
    .A2(_1114_),
    .B1(net25),
    .X(_1117_));
 sky130_fd_sc_hd__o211a_1 _1575_ (.A1(\product[28] ),
    .A2(_1114_),
    .B1(net25),
    .C1(\product[29] ),
    .X(_1118_));
 sky130_fd_sc_hd__o21ai_1 _1576_ (.A1(\product[29] ),
    .A2(_1117_),
    .B1(net136),
    .Y(_1119_));
 sky130_fd_sc_hd__a2bb2o_1 _1577_ (.A1_N(_1118_),
    .A2_N(_1119_),
    .B1(net87),
    .B2(net138),
    .X(_0124_));
 sky130_fd_sc_hd__o31a_1 _1578_ (.A1(\product[29] ),
    .A2(\product[28] ),
    .A3(_1114_),
    .B1(net25),
    .X(_1120_));
 sky130_fd_sc_hd__a21oi_1 _1579_ (.A1(\product[30] ),
    .A2(_1120_),
    .B1(_0870_),
    .Y(_1121_));
 sky130_fd_sc_hd__o21a_1 _1580_ (.A1(\product[30] ),
    .A2(_1120_),
    .B1(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__a31o_1 _1581_ (.A1(_0844_),
    .A2(net89),
    .A3(net142),
    .B1(_1122_),
    .X(_0125_));
 sky130_fd_sc_hd__or4_1 _1582_ (.A(\product[30] ),
    .B(\product[29] ),
    .C(\product[28] ),
    .D(_1114_),
    .X(_1123_));
 sky130_fd_sc_hd__a21oi_1 _1583_ (.A1(_1123_),
    .A2(net25),
    .B1(_0851_),
    .Y(_1124_));
 sky130_fd_sc_hd__a31o_1 _1584_ (.A1(_0851_),
    .A2(_1123_),
    .A3(net25),
    .B1(_0844_),
    .X(_1125_));
 sky130_fd_sc_hd__o221a_1 _1585_ (.A1(net139),
    .A2(net90),
    .B1(_1124_),
    .B2(_1125_),
    .C1(net142),
    .X(_0126_));
 sky130_fd_sc_hd__nor4_2 _1586_ (.A(\product[31] ),
    .B(\product[30] ),
    .C(\product[29] ),
    .D(\product[28] ),
    .Y(_1126_));
 sky130_fd_sc_hd__nand3b_4 _1587_ (.A_N(_1101_),
    .B(_1113_),
    .C(_1126_),
    .Y(_1127_));
 sky130_fd_sc_hd__a21oi_1 _1588_ (.A1(_1127_),
    .A2(net25),
    .B1(_0850_),
    .Y(_1128_));
 sky130_fd_sc_hd__a31o_1 _1589_ (.A1(_0850_),
    .A2(_1127_),
    .A3(net25),
    .B1(_0844_),
    .X(_1129_));
 sky130_fd_sc_hd__o221a_1 _1590_ (.A1(net139),
    .A2(net91),
    .B1(_1128_),
    .B2(_1129_),
    .C1(net142),
    .X(_0127_));
 sky130_fd_sc_hd__o21ai_1 _1591_ (.A1(\product[32] ),
    .A2(_1127_),
    .B1(net25),
    .Y(_1130_));
 sky130_fd_sc_hd__o21ai_1 _1592_ (.A1(\product[33] ),
    .A2(_1130_),
    .B1(net141),
    .Y(_1131_));
 sky130_fd_sc_hd__a21o_4 _1593_ (.A1(\product[33] ),
    .A2(_1130_),
    .B1(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__o211a_1 _1594_ (.A1(net141),
    .A2(net92),
    .B1(_0859_),
    .C1(_1132_),
    .X(_0128_));
 sky130_fd_sc_hd__or3_4 _1595_ (.A(\product[33] ),
    .B(\product[32] ),
    .C(_1127_),
    .X(_1133_));
 sky130_fd_sc_hd__a21oi_1 _1596_ (.A1(_1133_),
    .A2(net25),
    .B1(_0849_),
    .Y(_1134_));
 sky130_fd_sc_hd__a31o_1 _1597_ (.A1(_0849_),
    .A2(_1133_),
    .A3(net25),
    .B1(_0844_),
    .X(_1135_));
 sky130_fd_sc_hd__o221a_1 _1598_ (.A1(net141),
    .A2(net93),
    .B1(_1134_),
    .B2(_1135_),
    .C1(_0859_),
    .X(_0129_));
 sky130_fd_sc_hd__o21ai_1 _1599_ (.A1(\product[34] ),
    .A2(_1133_),
    .B1(net25),
    .Y(_1136_));
 sky130_fd_sc_hd__o21ai_1 _1600_ (.A1(\product[35] ),
    .A2(_1136_),
    .B1(net141),
    .Y(_1137_));
 sky130_fd_sc_hd__a21o_4 _1601_ (.A1(\product[35] ),
    .A2(_1136_),
    .B1(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__o211a_1 _1602_ (.A1(net141),
    .A2(net94),
    .B1(_0859_),
    .C1(_1138_),
    .X(_0130_));
 sky130_fd_sc_hd__o31ai_2 _1603_ (.A1(\product[35] ),
    .A2(\product[34] ),
    .A3(_1133_),
    .B1(net25),
    .Y(_1139_));
 sky130_fd_sc_hd__o21ai_1 _1604_ (.A1(\product[36] ),
    .A2(_1139_),
    .B1(net141),
    .Y(_1140_));
 sky130_fd_sc_hd__a21o_4 _1605_ (.A1(\product[36] ),
    .A2(_1139_),
    .B1(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__o211a_1 _1606_ (.A1(net141),
    .A2(net95),
    .B1(_0859_),
    .C1(_1141_),
    .X(_0131_));
 sky130_fd_sc_hd__o41ai_2 _1607_ (.A1(\product[36] ),
    .A2(\product[35] ),
    .A3(\product[34] ),
    .A4(_1133_),
    .B1(net25),
    .Y(_1142_));
 sky130_fd_sc_hd__o21ai_1 _1608_ (.A1(\product[37] ),
    .A2(_1142_),
    .B1(net141),
    .Y(_1143_));
 sky130_fd_sc_hd__a21o_4 _1609_ (.A1(\product[37] ),
    .A2(_1142_),
    .B1(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__o211a_1 _1610_ (.A1(net141),
    .A2(net96),
    .B1(_0859_),
    .C1(_1144_),
    .X(_0132_));
 sky130_fd_sc_hd__or4_1 _1611_ (.A(\product[37] ),
    .B(\product[36] ),
    .C(\product[35] ),
    .D(\product[34] ),
    .X(_1145_));
 sky130_fd_sc_hd__o21ai_2 _1612_ (.A1(_1133_),
    .A2(_1145_),
    .B1(net25),
    .Y(_1146_));
 sky130_fd_sc_hd__o21ai_1 _1613_ (.A1(\product[38] ),
    .A2(_1146_),
    .B1(net141),
    .Y(_1147_));
 sky130_fd_sc_hd__a21o_4 _1614_ (.A1(\product[38] ),
    .A2(_1146_),
    .B1(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__o211a_1 _1615_ (.A1(net141),
    .A2(net97),
    .B1(_0859_),
    .C1(_1148_),
    .X(_0133_));
 sky130_fd_sc_hd__nand2_1 _1616_ (.A(\product[38] ),
    .B(net25),
    .Y(_1149_));
 sky130_fd_sc_hd__a21oi_1 _1617_ (.A1(_1146_),
    .A2(_1149_),
    .B1(\product[39] ),
    .Y(_1150_));
 sky130_fd_sc_hd__a31o_1 _1618_ (.A1(\product[39] ),
    .A2(_1146_),
    .A3(_1149_),
    .B1(_0844_),
    .X(_1151_));
 sky130_fd_sc_hd__o221a_1 _1619_ (.A1(net141),
    .A2(net98),
    .B1(_1150_),
    .B2(_1151_),
    .C1(_0859_),
    .X(_0134_));
 sky130_fd_sc_hd__or3_1 _1620_ (.A(\product[39] ),
    .B(\product[33] ),
    .C(\product[32] ),
    .X(_1152_));
 sky130_fd_sc_hd__nor3_2 _1621_ (.A(_1152_),
    .B(\product[38] ),
    .C(_1145_),
    .Y(_1153_));
 sky130_fd_sc_hd__nand4b_4 _1622_ (.A_N(_1101_),
    .B(_1113_),
    .C(_1126_),
    .D(net134),
    .Y(_1154_));
 sky130_fd_sc_hd__a21oi_1 _1623_ (.A1(_1154_),
    .A2(net25),
    .B1(_0848_),
    .Y(_1155_));
 sky130_fd_sc_hd__a31o_1 _1624_ (.A1(_0848_),
    .A2(_1154_),
    .A3(net25),
    .B1(_0844_),
    .X(_1156_));
 sky130_fd_sc_hd__o221a_1 _1625_ (.A1(net139),
    .A2(net100),
    .B1(_1155_),
    .B2(_1156_),
    .C1(net142),
    .X(_0135_));
 sky130_fd_sc_hd__o21ai_1 _1626_ (.A1(\product[40] ),
    .A2(_1154_),
    .B1(net25),
    .Y(_1157_));
 sky130_fd_sc_hd__o21ai_1 _1627_ (.A1(\product[41] ),
    .A2(_1157_),
    .B1(net140),
    .Y(_1158_));
 sky130_fd_sc_hd__a21o_4 _1628_ (.A1(\product[41] ),
    .A2(_1157_),
    .B1(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__o211a_1 _1629_ (.A1(net139),
    .A2(net101),
    .B1(net142),
    .C1(_1159_),
    .X(_0136_));
 sky130_fd_sc_hd__o31ai_2 _1630_ (.A1(\product[41] ),
    .A2(\product[40] ),
    .A3(_1154_),
    .B1(net25),
    .Y(_1160_));
 sky130_fd_sc_hd__o21ai_1 _1631_ (.A1(\product[42] ),
    .A2(_1160_),
    .B1(net140),
    .Y(_1161_));
 sky130_fd_sc_hd__a21o_4 _1632_ (.A1(\product[42] ),
    .A2(_1160_),
    .B1(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__o211a_1 _1633_ (.A1(net139),
    .A2(net102),
    .B1(net142),
    .C1(_1162_),
    .X(_0137_));
 sky130_fd_sc_hd__or4_4 _1634_ (.A(\product[42] ),
    .B(\product[41] ),
    .C(\product[40] ),
    .D(_1154_),
    .X(_1163_));
 sky130_fd_sc_hd__nand2_1 _1635_ (.A(_1163_),
    .B(net25),
    .Y(_1164_));
 sky130_fd_sc_hd__nor2_1 _1636_ (.A(\product[43] ),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__a21o_1 _1637_ (.A1(_1164_),
    .A2(\product[43] ),
    .B1(_0844_),
    .X(_1166_));
 sky130_fd_sc_hd__o221a_1 _1638_ (.A1(net140),
    .A2(net103),
    .B1(_1165_),
    .B2(_1166_),
    .C1(_0859_),
    .X(_0138_));
 sky130_fd_sc_hd__nor4_4 _1639_ (.A(\product[43] ),
    .B(\product[42] ),
    .C(\product[41] ),
    .D(\product[40] ),
    .Y(_1167_));
 sky130_fd_sc_hd__nand3b_4 _1640_ (.A_N(_1127_),
    .B(_1153_),
    .C(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__a21oi_1 _1641_ (.A1(_1168_),
    .A2(net25),
    .B1(_0847_),
    .Y(_1169_));
 sky130_fd_sc_hd__a31o_1 _1642_ (.A1(_0847_),
    .A2(_1168_),
    .A3(net25),
    .B1(_0844_),
    .X(_1170_));
 sky130_fd_sc_hd__o221a_1 _1643_ (.A1(net140),
    .A2(net104),
    .B1(_1169_),
    .B2(_1170_),
    .C1(_0859_),
    .X(_0139_));
 sky130_fd_sc_hd__o31a_1 _1644_ (.A1(\product[44] ),
    .A2(\product[43] ),
    .A3(_1163_),
    .B1(net25),
    .X(_1171_));
 sky130_fd_sc_hd__o311a_1 _1645_ (.A1(\product[44] ),
    .A2(\product[43] ),
    .A3(_1163_),
    .B1(net25),
    .C1(\product[45] ),
    .X(_1172_));
 sky130_fd_sc_hd__o21ai_1 _1646_ (.A1(\product[45] ),
    .A2(_1171_),
    .B1(net135),
    .Y(_1173_));
 sky130_fd_sc_hd__a2bb2o_1 _1647_ (.A1_N(_1172_),
    .A2_N(_1173_),
    .B1(net105),
    .B2(net137),
    .X(_0140_));
 sky130_fd_sc_hd__or4_1 _1648_ (.A(\product[45] ),
    .B(\product[44] ),
    .C(\product[43] ),
    .D(_1163_),
    .X(_1174_));
 sky130_fd_sc_hd__o31a_1 _1649_ (.A1(\product[45] ),
    .A2(\product[44] ),
    .A3(_1168_),
    .B1(net25),
    .X(_1175_));
 sky130_fd_sc_hd__a21oi_1 _1650_ (.A1(_1174_),
    .A2(net25),
    .B1(_0846_),
    .Y(_1176_));
 sky130_fd_sc_hd__a31o_1 _1651_ (.A1(_0846_),
    .A2(_1174_),
    .A3(net25),
    .B1(_0844_),
    .X(_0230_));
 sky130_fd_sc_hd__o221a_1 _1652_ (.A1(net140),
    .A2(net106),
    .B1(_0230_),
    .B2(_1176_),
    .C1(_0859_),
    .X(_0141_));
 sky130_fd_sc_hd__a211o_1 _1653_ (.A1(\product[46] ),
    .A2(net25),
    .B1(_1175_),
    .C1(\product[47] ),
    .X(_0231_));
 sky130_fd_sc_hd__o211ai_1 _1654_ (.A1(\product[46] ),
    .A2(_1174_),
    .B1(net25),
    .C1(\product[47] ),
    .Y(_0232_));
 sky130_fd_sc_hd__a32o_1 _1655_ (.A1(_0232_),
    .A2(net135),
    .A3(_0231_),
    .B1(net137),
    .B2(net107),
    .X(_0142_));
 sky130_fd_sc_hd__nor4_2 _1656_ (.A(\product[47] ),
    .B(\product[46] ),
    .C(\product[45] ),
    .D(\product[44] ),
    .Y(_0233_));
 sky130_fd_sc_hd__nand3b_4 _1657_ (.A_N(_1154_),
    .B(_1167_),
    .C(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__a21oi_1 _1658_ (.A1(_0234_),
    .A2(net25),
    .B1(_0845_),
    .Y(_0235_));
 sky130_fd_sc_hd__a31o_1 _1659_ (.A1(_0845_),
    .A2(_0234_),
    .A3(net25),
    .B1(_0844_),
    .X(_0236_));
 sky130_fd_sc_hd__o221a_1 _1660_ (.A1(net141),
    .A2(net108),
    .B1(_0235_),
    .B2(_0236_),
    .C1(_0859_),
    .X(_0143_));
 sky130_fd_sc_hd__o21ai_1 _1661_ (.A1(\product[48] ),
    .A2(_0234_),
    .B1(net25),
    .Y(_0237_));
 sky130_fd_sc_hd__o21ai_1 _1662_ (.A1(\product[49] ),
    .A2(_0237_),
    .B1(net140),
    .Y(_0238_));
 sky130_fd_sc_hd__a21o_4 _1663_ (.A1(\product[49] ),
    .A2(_0237_),
    .B1(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__o211a_1 _1664_ (.A1(net140),
    .A2(net109),
    .B1(_0859_),
    .C1(_0239_),
    .X(_0144_));
 sky130_fd_sc_hd__or2_4 _1665_ (.A(\product[49] ),
    .B(\product[48] ),
    .X(_0240_));
 sky130_fd_sc_hd__o31a_1 _1666_ (.A1(\product[49] ),
    .A2(\product[48] ),
    .A3(_0234_),
    .B1(net25),
    .X(_0241_));
 sky130_fd_sc_hd__o21ai_2 _1667_ (.A1(_0234_),
    .A2(_0240_),
    .B1(net25),
    .Y(_0242_));
 sky130_fd_sc_hd__o21ai_1 _1668_ (.A1(\product[50] ),
    .A2(_0242_),
    .B1(net141),
    .Y(_0243_));
 sky130_fd_sc_hd__a21o_4 _1669_ (.A1(\product[50] ),
    .A2(_0242_),
    .B1(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__o211a_1 _1670_ (.A1(net141),
    .A2(net111),
    .B1(_0859_),
    .C1(_0244_),
    .X(_0145_));
 sky130_fd_sc_hd__nand2_1 _1671_ (.A(\product[50] ),
    .B(net25),
    .Y(_0245_));
 sky130_fd_sc_hd__a21oi_1 _1672_ (.A1(_0242_),
    .A2(_0245_),
    .B1(\product[51] ),
    .Y(_0246_));
 sky130_fd_sc_hd__a31o_1 _1673_ (.A1(_0242_),
    .A2(_0245_),
    .A3(\product[51] ),
    .B1(_0844_),
    .X(_0247_));
 sky130_fd_sc_hd__o221a_1 _1674_ (.A1(net141),
    .A2(net112),
    .B1(_0246_),
    .B2(_0247_),
    .C1(_0859_),
    .X(_0146_));
 sky130_fd_sc_hd__o41ai_4 _1675_ (.A1(\product[51] ),
    .A2(_0240_),
    .A3(\product[50] ),
    .A4(_0234_),
    .B1(net25),
    .Y(_0248_));
 sky130_fd_sc_hd__o21ai_1 _1676_ (.A1(\product[52] ),
    .A2(_0248_),
    .B1(net141),
    .Y(_0249_));
 sky130_fd_sc_hd__a21o_4 _1677_ (.A1(\product[52] ),
    .A2(_0248_),
    .B1(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__o211a_1 _1678_ (.A1(net141),
    .A2(net113),
    .B1(_0859_),
    .C1(_0250_),
    .X(_0147_));
 sky130_fd_sc_hd__nand2_1 _1679_ (.A(\product[52] ),
    .B(net25),
    .Y(_0251_));
 sky130_fd_sc_hd__a21oi_1 _1680_ (.A1(_0248_),
    .A2(_0251_),
    .B1(\product[53] ),
    .Y(_0252_));
 sky130_fd_sc_hd__a31o_1 _1681_ (.A1(_0248_),
    .A2(_0251_),
    .A3(\product[53] ),
    .B1(_0844_),
    .X(_0253_));
 sky130_fd_sc_hd__o221a_1 _1682_ (.A1(net141),
    .A2(net114),
    .B1(_0252_),
    .B2(_0253_),
    .C1(_0859_),
    .X(_0148_));
 sky130_fd_sc_hd__or4_4 _1683_ (.A(\product[53] ),
    .B(\product[52] ),
    .C(\product[51] ),
    .D(\product[50] ),
    .X(_0254_));
 sky130_fd_sc_hd__a211o_1 _1684_ (.A1(_0254_),
    .A2(net25),
    .B1(\product[54] ),
    .C1(_0241_),
    .X(_0255_));
 sky130_fd_sc_hd__o311ai_2 _1685_ (.A1(_0234_),
    .A2(_0240_),
    .A3(_0254_),
    .B1(net25),
    .C1(\product[54] ),
    .Y(_0256_));
 sky130_fd_sc_hd__a32o_1 _1686_ (.A1(_0255_),
    .A2(_0256_),
    .A3(net135),
    .B1(net137),
    .B2(net115),
    .X(_0149_));
 sky130_fd_sc_hd__o31a_1 _1687_ (.A1(\product[54] ),
    .A2(_0254_),
    .A3(_0241_),
    .B1(net25),
    .X(_0257_));
 sky130_fd_sc_hd__xor2_4 _1688_ (.A(\product[55] ),
    .B(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__a22o_1 _1689_ (.A1(net116),
    .A2(net137),
    .B1(_0258_),
    .B2(net135),
    .X(_0150_));
 sky130_fd_sc_hd__or4_4 _1690_ (.A(\product[55] ),
    .B(\product[54] ),
    .C(_0240_),
    .D(_0254_),
    .X(_0259_));
 sky130_fd_sc_hd__or2_2 _1691_ (.A(_0234_),
    .B(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__o21ai_1 _1692_ (.A1(_0234_),
    .A2(_0259_),
    .B1(net25),
    .Y(_0261_));
 sky130_fd_sc_hd__o21ai_1 _1693_ (.A1(\product[56] ),
    .A2(_0261_),
    .B1(net140),
    .Y(_0262_));
 sky130_fd_sc_hd__a21o_1 _1694_ (.A1(\product[56] ),
    .A2(_0261_),
    .B1(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__o211a_1 _1695_ (.A1(net140),
    .A2(net117),
    .B1(_0859_),
    .C1(_0263_),
    .X(_0151_));
 sky130_fd_sc_hd__o21ai_1 _1696_ (.A1(\product[56] ),
    .A2(_0260_),
    .B1(net25),
    .Y(_0264_));
 sky130_fd_sc_hd__o21ai_1 _1697_ (.A1(\product[57] ),
    .A2(_0264_),
    .B1(net140),
    .Y(_0265_));
 sky130_fd_sc_hd__a21o_1 _1698_ (.A1(\product[57] ),
    .A2(_0264_),
    .B1(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__o211a_1 _1699_ (.A1(net140),
    .A2(net118),
    .B1(_0859_),
    .C1(_0266_),
    .X(_0152_));
 sky130_fd_sc_hd__o31ai_1 _1700_ (.A1(\product[57] ),
    .A2(\product[56] ),
    .A3(_0260_),
    .B1(net25),
    .Y(_0267_));
 sky130_fd_sc_hd__o21ai_1 _1701_ (.A1(\product[58] ),
    .A2(_0267_),
    .B1(net140),
    .Y(_0268_));
 sky130_fd_sc_hd__a21o_1 _1702_ (.A1(\product[58] ),
    .A2(_0267_),
    .B1(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__o211a_1 _1703_ (.A1(net140),
    .A2(net119),
    .B1(_0859_),
    .C1(_0269_),
    .X(_0153_));
 sky130_fd_sc_hd__o41ai_1 _1704_ (.A1(\product[58] ),
    .A2(\product[57] ),
    .A3(\product[56] ),
    .A4(_0260_),
    .B1(net25),
    .Y(_0270_));
 sky130_fd_sc_hd__nand2_1 _1705_ (.A(\product[59] ),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__o21a_1 _1706_ (.A1(\product[59] ),
    .A2(_0270_),
    .B1(net140),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_1 _1707_ (.A(_0272_),
    .B(_0271_),
    .Y(_0273_));
 sky130_fd_sc_hd__o211a_1 _1708_ (.A1(net140),
    .A2(net120),
    .B1(_0859_),
    .C1(_0273_),
    .X(_0154_));
 sky130_fd_sc_hd__or4_1 _1709_ (.A(\product[59] ),
    .B(\product[58] ),
    .C(\product[57] ),
    .D(\product[56] ),
    .X(_0274_));
 sky130_fd_sc_hd__o21ai_4 _1710_ (.A1(_0260_),
    .A2(_0274_),
    .B1(net25),
    .Y(_0275_));
 sky130_fd_sc_hd__o21ai_1 _1711_ (.A1(\product[60] ),
    .A2(_0275_),
    .B1(net140),
    .Y(_0276_));
 sky130_fd_sc_hd__a21o_1 _1712_ (.A1(\product[60] ),
    .A2(_0275_),
    .B1(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__o211a_1 _1713_ (.A1(net140),
    .A2(net122),
    .B1(_0859_),
    .C1(_0277_),
    .X(_0155_));
 sky130_fd_sc_hd__nand2_1 _1714_ (.A(\product[60] ),
    .B(net25),
    .Y(_0278_));
 sky130_fd_sc_hd__a21oi_1 _1715_ (.A1(_0275_),
    .A2(_0278_),
    .B1(\product[61] ),
    .Y(_0279_));
 sky130_fd_sc_hd__a31o_1 _1716_ (.A1(_0275_),
    .A2(_0278_),
    .A3(\product[61] ),
    .B1(_0844_),
    .X(_0280_));
 sky130_fd_sc_hd__o221a_1 _1717_ (.A1(net140),
    .A2(net123),
    .B1(_0279_),
    .B2(_0280_),
    .C1(_0859_),
    .X(_0156_));
 sky130_fd_sc_hd__o21ai_2 _1718_ (.A1(\product[61] ),
    .A2(\product[60] ),
    .B1(net25),
    .Y(_0281_));
 sky130_fd_sc_hd__a21oi_1 _1719_ (.A1(_0275_),
    .A2(_0281_),
    .B1(\product[62] ),
    .Y(_0282_));
 sky130_fd_sc_hd__a31o_1 _1720_ (.A1(_0275_),
    .A2(_0281_),
    .A3(\product[62] ),
    .B1(_0844_),
    .X(_0283_));
 sky130_fd_sc_hd__o221a_1 _1721_ (.A1(net140),
    .A2(net124),
    .B1(_0282_),
    .B2(_0283_),
    .C1(_0859_),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_1 _1722_ (.A(\product[62] ),
    .B(net25),
    .Y(_0284_));
 sky130_fd_sc_hd__a31oi_1 _1723_ (.A1(_0275_),
    .A2(_0281_),
    .A3(_0284_),
    .B1(\product[63] ),
    .Y(_0285_));
 sky130_fd_sc_hd__a41o_1 _1724_ (.A1(_0275_),
    .A2(_0281_),
    .A3(_0284_),
    .A4(\product[63] ),
    .B1(_0844_),
    .X(_0286_));
 sky130_fd_sc_hd__o221a_1 _1725_ (.A1(net140),
    .A2(net125),
    .B1(_0285_),
    .B2(_0286_),
    .C1(_0859_),
    .X(_0158_));
 sky130_fd_sc_hd__and2_4 _1726_ (.A(_0844_),
    .B(\multiplier[0] ),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_8 _1727_ (.A(_0844_),
    .B(\multiplier[0] ),
    .Y(_0288_));
 sky130_fd_sc_hd__a21oi_1 _1728_ (.A1(\multiplicand[0] ),
    .A2(net133),
    .B1(\product[0] ),
    .Y(_0289_));
 sky130_fd_sc_hd__a311oi_1 _1729_ (.A1(\product[0] ),
    .A2(\multiplicand[0] ),
    .A3(net133),
    .B1(_0289_),
    .C1(net65),
    .Y(_0159_));
 sky130_fd_sc_hd__a21o_1 _1730_ (.A1(\product[0] ),
    .A2(\multiplicand[0] ),
    .B1(\multiplicand[1] ),
    .X(_0290_));
 sky130_fd_sc_hd__nand3_1 _1731_ (.A(\product[0] ),
    .B(\multiplicand[0] ),
    .C(\multiplicand[1] ),
    .Y(_0291_));
 sky130_fd_sc_hd__a31o_1 _1732_ (.A1(net133),
    .A2(_0290_),
    .A3(_0291_),
    .B1(\product[1] ),
    .X(_0292_));
 sky130_fd_sc_hd__nand4_1 _1733_ (.A(\product[1] ),
    .B(net133),
    .C(_0290_),
    .D(_0291_),
    .Y(_0293_));
 sky130_fd_sc_hd__and2_1 _1734_ (.A(\product[1] ),
    .B(\multiplicand[1] ),
    .X(_0294_));
 sky130_fd_sc_hd__o211a_1 _1735_ (.A1(\product[1] ),
    .A2(\multiplicand[1] ),
    .B1(\multiplicand[0] ),
    .C1(\product[0] ),
    .X(_0295_));
 sky130_fd_sc_hd__and3_1 _1736_ (.A(net142),
    .B(_0292_),
    .C(_0293_),
    .X(_0160_));
 sky130_fd_sc_hd__nand2_1 _1737_ (.A(\product[2] ),
    .B(\multiplicand[2] ),
    .Y(_0296_));
 sky130_fd_sc_hd__or2_1 _1738_ (.A(\product[2] ),
    .B(\multiplicand[2] ),
    .X(_0297_));
 sky130_fd_sc_hd__and2b_1 _1739_ (.A_N(\product[2] ),
    .B(\multiplicand[2] ),
    .X(_0298_));
 sky130_fd_sc_hd__and2b_1 _1740_ (.A_N(\multiplicand[2] ),
    .B(\product[2] ),
    .X(_0299_));
 sky130_fd_sc_hd__a22o_1 _1741_ (.A1(\product[0] ),
    .A2(\multiplicand[0] ),
    .B1(\multiplicand[1] ),
    .B2(\product[1] ),
    .X(_0300_));
 sky130_fd_sc_hd__or4_1 _1742_ (.A(_0294_),
    .B(_0295_),
    .C(_0298_),
    .D(_0299_),
    .X(_0301_));
 sky130_fd_sc_hd__o2111ai_4 _1743_ (.A1(\product[1] ),
    .A2(\multiplicand[1] ),
    .B1(_0296_),
    .C1(_0297_),
    .D1(_0300_),
    .Y(_0302_));
 sky130_fd_sc_hd__a21o_1 _1744_ (.A1(_0301_),
    .A2(_0302_),
    .B1(net131),
    .X(_0303_));
 sky130_fd_sc_hd__o211a_1 _1745_ (.A1(\product[2] ),
    .A2(net133),
    .B1(_0303_),
    .C1(net142),
    .X(_0161_));
 sky130_fd_sc_hd__nor2_1 _1746_ (.A(\product[3] ),
    .B(\multiplicand[3] ),
    .Y(_0304_));
 sky130_fd_sc_hd__or2_4 _1747_ (.A(\product[3] ),
    .B(\multiplicand[3] ),
    .X(_0305_));
 sky130_fd_sc_hd__and2_1 _1748_ (.A(\product[3] ),
    .B(\multiplicand[3] ),
    .X(_0306_));
 sky130_fd_sc_hd__nor2_1 _1749_ (.A(_0304_),
    .B(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__o2bb2a_1 _1750_ (.A1_N(_0296_),
    .A2_N(_0302_),
    .B1(_0304_),
    .B2(_0306_),
    .X(_0308_));
 sky130_fd_sc_hd__a21oi_1 _1751_ (.A1(\product[2] ),
    .A2(\multiplicand[2] ),
    .B1(_0306_),
    .Y(_0309_));
 sky130_fd_sc_hd__nand2_2 _1752_ (.A(_0302_),
    .B(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__a31o_1 _1753_ (.A1(_0302_),
    .A2(_0305_),
    .A3(_0309_),
    .B1(net131),
    .X(_0311_));
 sky130_fd_sc_hd__o221a_1 _1754_ (.A1(\product[3] ),
    .A2(net133),
    .B1(_0311_),
    .B2(_0308_),
    .C1(net142),
    .X(_0162_));
 sky130_fd_sc_hd__nor2_1 _1755_ (.A(\product[4] ),
    .B(\multiplicand[4] ),
    .Y(_0312_));
 sky130_fd_sc_hd__and2_1 _1756_ (.A(\product[4] ),
    .B(\multiplicand[4] ),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _1757_ (.A(\product[4] ),
    .B(\multiplicand[4] ),
    .Y(_0314_));
 sky130_fd_sc_hd__nor2_1 _1758_ (.A(_0312_),
    .B(_0313_),
    .Y(_0315_));
 sky130_fd_sc_hd__o221ai_4 _1759_ (.A1(_0294_),
    .A2(_0295_),
    .B1(_0298_),
    .B2(_0299_),
    .C1(_0307_),
    .Y(_0316_));
 sky130_fd_sc_hd__a31oi_2 _1760_ (.A1(_0305_),
    .A2(\multiplicand[2] ),
    .A3(\product[2] ),
    .B1(_0306_),
    .Y(_0317_));
 sky130_fd_sc_hd__o31a_1 _1761_ (.A1(_0304_),
    .A2(_0306_),
    .A3(_0302_),
    .B1(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__or3_1 _1762_ (.A(_0312_),
    .B(_0313_),
    .C(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__a21o_1 _1763_ (.A1(_0305_),
    .A2(_0310_),
    .B1(_0315_),
    .X(_0320_));
 sky130_fd_sc_hd__a21o_1 _1764_ (.A1(_0319_),
    .A2(_0320_),
    .B1(net131),
    .X(_0321_));
 sky130_fd_sc_hd__o211a_1 _1765_ (.A1(\product[4] ),
    .A2(net133),
    .B1(_0321_),
    .C1(net142),
    .X(_0163_));
 sky130_fd_sc_hd__nor2_2 _1766_ (.A(\product[5] ),
    .B(\multiplicand[5] ),
    .Y(_0322_));
 sky130_fd_sc_hd__and2_1 _1767_ (.A(\product[5] ),
    .B(\multiplicand[5] ),
    .X(_0323_));
 sky130_fd_sc_hd__nand2_1 _1768_ (.A(\product[5] ),
    .B(\multiplicand[5] ),
    .Y(_0324_));
 sky130_fd_sc_hd__nor2_1 _1769_ (.A(_0322_),
    .B(_0323_),
    .Y(_0325_));
 sky130_fd_sc_hd__o2bb2a_1 _1770_ (.A1_N(_0314_),
    .A2_N(_0319_),
    .B1(_0322_),
    .B2(_0323_),
    .X(_0326_));
 sky130_fd_sc_hd__a31o_1 _1771_ (.A1(_0314_),
    .A2(_0319_),
    .A3(_0325_),
    .B1(net131),
    .X(_0327_));
 sky130_fd_sc_hd__o221a_1 _1772_ (.A1(\product[5] ),
    .A2(net133),
    .B1(_0327_),
    .B2(_0326_),
    .C1(net142),
    .X(_0164_));
 sky130_fd_sc_hd__nor2_1 _1773_ (.A(\product[6] ),
    .B(\multiplicand[6] ),
    .Y(_0328_));
 sky130_fd_sc_hd__or2_1 _1774_ (.A(\product[6] ),
    .B(\multiplicand[6] ),
    .X(_0329_));
 sky130_fd_sc_hd__and2_1 _1775_ (.A(\product[6] ),
    .B(\multiplicand[6] ),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _1776_ (.A(\product[6] ),
    .B(\multiplicand[6] ),
    .Y(_0331_));
 sky130_fd_sc_hd__nor2_1 _1777_ (.A(_0328_),
    .B(_0330_),
    .Y(_0332_));
 sky130_fd_sc_hd__o21a_1 _1778_ (.A1(_0314_),
    .A2(_0322_),
    .B1(_0324_),
    .X(_0333_));
 sky130_fd_sc_hd__o21ai_1 _1779_ (.A1(_0314_),
    .A2(_0322_),
    .B1(_0324_),
    .Y(_0334_));
 sky130_fd_sc_hd__nor4_2 _1780_ (.A(_0312_),
    .B(_0313_),
    .C(_0322_),
    .D(_0323_),
    .Y(_0335_));
 sky130_fd_sc_hd__or4b_1 _1781_ (.A(_0312_),
    .B(_0313_),
    .C(_0318_),
    .D_N(_0325_),
    .X(_0336_));
 sky130_fd_sc_hd__or3b_1 _1782_ (.A(_0332_),
    .B(_0334_),
    .C_N(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__a211o_1 _1783_ (.A1(_0336_),
    .A2(_0333_),
    .B1(_0330_),
    .C1(_0328_),
    .X(_0338_));
 sky130_fd_sc_hd__a21o_1 _1784_ (.A1(_0337_),
    .A2(_0338_),
    .B1(net131),
    .X(_0339_));
 sky130_fd_sc_hd__o211a_1 _1785_ (.A1(\product[6] ),
    .A2(net133),
    .B1(_0339_),
    .C1(net142),
    .X(_0165_));
 sky130_fd_sc_hd__nor2_1 _1786_ (.A(\product[7] ),
    .B(\multiplicand[7] ),
    .Y(_0340_));
 sky130_fd_sc_hd__and2_1 _1787_ (.A(\product[7] ),
    .B(\multiplicand[7] ),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_2 _1788_ (.A(_0340_),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__o2bb2a_1 _1789_ (.A1_N(_0331_),
    .A2_N(_0338_),
    .B1(_0340_),
    .B2(_0341_),
    .X(_0343_));
 sky130_fd_sc_hd__a31o_1 _1790_ (.A1(_0331_),
    .A2(_0338_),
    .A3(_0342_),
    .B1(net131),
    .X(_0344_));
 sky130_fd_sc_hd__o221a_1 _1791_ (.A1(\product[7] ),
    .A2(net133),
    .B1(_0344_),
    .B2(_0343_),
    .C1(net142),
    .X(_0166_));
 sky130_fd_sc_hd__and3_1 _1792_ (.A(_0342_),
    .B(_0331_),
    .C(_0329_),
    .X(_0345_));
 sky130_fd_sc_hd__nand4_2 _1793_ (.A(_0315_),
    .B(_0325_),
    .C(_0332_),
    .D(_0342_),
    .Y(_0346_));
 sky130_fd_sc_hd__a21oi_4 _1794_ (.A1(_0316_),
    .A2(_0317_),
    .B1(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__o21bai_1 _1795_ (.A1(_0331_),
    .A2(_0340_),
    .B1_N(_0341_),
    .Y(_0348_));
 sky130_fd_sc_hd__a31o_4 _1796_ (.A1(_0332_),
    .A2(_0342_),
    .A3(_0334_),
    .B1(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__a41oi_4 _1797_ (.A1(_0345_),
    .A2(_0310_),
    .A3(_0305_),
    .A4(_0335_),
    .B1(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__a41o_4 _1798_ (.A1(_0345_),
    .A2(_0310_),
    .A3(_0305_),
    .A4(_0335_),
    .B1(_0349_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _1799_ (.A(\product[8] ),
    .B(\multiplicand[8] ),
    .Y(_0352_));
 sky130_fd_sc_hd__or2_1 _1800_ (.A(\product[8] ),
    .B(\multiplicand[8] ),
    .X(_0353_));
 sky130_fd_sc_hd__a21oi_1 _1801_ (.A1(_0352_),
    .A2(_0353_),
    .B1(_0351_),
    .Y(_0354_));
 sky130_fd_sc_hd__and3_1 _1802_ (.A(_0351_),
    .B(_0352_),
    .C(_0353_),
    .X(_0355_));
 sky130_fd_sc_hd__o21ai_1 _1803_ (.A1(_0354_),
    .A2(_0355_),
    .B1(net132),
    .Y(_0356_));
 sky130_fd_sc_hd__o211a_1 _1804_ (.A1(\product[8] ),
    .A2(net132),
    .B1(_0356_),
    .C1(net142),
    .X(_0167_));
 sky130_fd_sc_hd__a21oi_1 _1805_ (.A1(\product[8] ),
    .A2(\multiplicand[8] ),
    .B1(_0355_),
    .Y(_0357_));
 sky130_fd_sc_hd__or2_2 _1806_ (.A(\product[9] ),
    .B(\multiplicand[9] ),
    .X(_0358_));
 sky130_fd_sc_hd__nand2_1 _1807_ (.A(\product[9] ),
    .B(\multiplicand[9] ),
    .Y(_0359_));
 sky130_fd_sc_hd__and2b_1 _1808_ (.A_N(\product[9] ),
    .B(\multiplicand[9] ),
    .X(_0360_));
 sky130_fd_sc_hd__nor2_1 _1809_ (.A(\multiplicand[9] ),
    .B(_0856_),
    .Y(_0361_));
 sky130_fd_sc_hd__or3_1 _1810_ (.A(_0357_),
    .B(_0360_),
    .C(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__a31oi_1 _1811_ (.A1(_0357_),
    .A2(_0358_),
    .A3(_0359_),
    .B1(net131),
    .Y(_0363_));
 sky130_fd_sc_hd__a221oi_1 _1812_ (.A1(_0856_),
    .A2(net131),
    .B1(_0362_),
    .B2(_0363_),
    .C1(net65),
    .Y(_0168_));
 sky130_fd_sc_hd__nand2b_1 _1813_ (.A_N(\product[10] ),
    .B(\multiplicand[10] ),
    .Y(_0364_));
 sky130_fd_sc_hd__nand2b_1 _1814_ (.A_N(\multiplicand[10] ),
    .B(\product[10] ),
    .Y(_0365_));
 sky130_fd_sc_hd__nand2_2 _1815_ (.A(_0364_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__o21ai_1 _1816_ (.A1(\product[9] ),
    .A2(\multiplicand[9] ),
    .B1(\multiplicand[8] ),
    .Y(_0367_));
 sky130_fd_sc_hd__o21ai_2 _1817_ (.A1(_0857_),
    .A2(_0367_),
    .B1(_0359_),
    .Y(_0368_));
 sky130_fd_sc_hd__a221o_1 _1818_ (.A1(\product[8] ),
    .A2(\multiplicand[8] ),
    .B1(\multiplicand[9] ),
    .B2(\product[9] ),
    .C1(_0355_),
    .X(_0369_));
 sky130_fd_sc_hd__nand4_2 _1819_ (.A(_0352_),
    .B(_0353_),
    .C(_0358_),
    .D(_0359_),
    .Y(_0370_));
 sky130_fd_sc_hd__a211o_1 _1820_ (.A1(_0355_),
    .A2(_0358_),
    .B1(_0366_),
    .C1(_0368_),
    .X(_0371_));
 sky130_fd_sc_hd__o211ai_1 _1821_ (.A1(\product[9] ),
    .A2(\multiplicand[9] ),
    .B1(_0366_),
    .C1(_0369_),
    .Y(_0372_));
 sky130_fd_sc_hd__a21o_1 _1822_ (.A1(_0371_),
    .A2(_0372_),
    .B1(net131),
    .X(_0373_));
 sky130_fd_sc_hd__o211a_1 _1823_ (.A1(\product[10] ),
    .A2(net132),
    .B1(_0373_),
    .C1(net142),
    .X(_0169_));
 sky130_fd_sc_hd__a32oi_2 _1824_ (.A1(_0358_),
    .A2(_0369_),
    .A3(_0366_),
    .B1(\product[10] ),
    .B2(\multiplicand[10] ),
    .Y(_0374_));
 sky130_fd_sc_hd__nand2b_1 _1825_ (.A_N(\product[11] ),
    .B(\multiplicand[11] ),
    .Y(_0375_));
 sky130_fd_sc_hd__nand2b_1 _1826_ (.A_N(\multiplicand[11] ),
    .B(\product[11] ),
    .Y(_0376_));
 sky130_fd_sc_hd__nand2_2 _1827_ (.A(_0375_),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__o21ai_1 _1828_ (.A1(_0374_),
    .A2(_0377_),
    .B1(net132),
    .Y(_0378_));
 sky130_fd_sc_hd__a21o_1 _1829_ (.A1(_0374_),
    .A2(_0377_),
    .B1(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__o211a_1 _1830_ (.A1(\product[11] ),
    .A2(net132),
    .B1(_0379_),
    .C1(net142),
    .X(_0170_));
 sky130_fd_sc_hd__a22o_1 _1831_ (.A1(_0364_),
    .A2(_0365_),
    .B1(_0375_),
    .B2(_0376_),
    .X(_0380_));
 sky130_fd_sc_hd__o21a_1 _1832_ (.A1(\product[11] ),
    .A2(\multiplicand[11] ),
    .B1(\multiplicand[10] ),
    .X(_0381_));
 sky130_fd_sc_hd__a22o_1 _1833_ (.A1(\product[11] ),
    .A2(\multiplicand[11] ),
    .B1(_0381_),
    .B2(\product[10] ),
    .X(_0382_));
 sky130_fd_sc_hd__a31oi_4 _1834_ (.A1(_0366_),
    .A2(_0368_),
    .A3(_0377_),
    .B1(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__o211a_1 _1835_ (.A1(_0360_),
    .A2(_0361_),
    .B1(_0366_),
    .C1(_0377_),
    .X(_0384_));
 sky130_fd_sc_hd__or3_1 _1836_ (.A(_0370_),
    .B(_0380_),
    .C(net130),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _1837_ (.A(\product[12] ),
    .B(\multiplicand[12] ),
    .X(_0386_));
 sky130_fd_sc_hd__nor2_1 _1838_ (.A(\product[12] ),
    .B(\multiplicand[12] ),
    .Y(_0387_));
 sky130_fd_sc_hd__nor2_1 _1839_ (.A(_0386_),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__or2_1 _1840_ (.A(_0386_),
    .B(_0387_),
    .X(_0389_));
 sky130_fd_sc_hd__o311a_1 _1841_ (.A1(_0370_),
    .A2(_0380_),
    .A3(net130),
    .B1(_0383_),
    .C1(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__a21oi_4 _1842_ (.A1(_0385_),
    .A2(_0383_),
    .B1(_0389_),
    .Y(_0391_));
 sky130_fd_sc_hd__o21ai_1 _1843_ (.A1(_0390_),
    .A2(_0391_),
    .B1(net132),
    .Y(_0392_));
 sky130_fd_sc_hd__o211a_1 _1844_ (.A1(\product[12] ),
    .A2(net132),
    .B1(_0392_),
    .C1(net142),
    .X(_0171_));
 sky130_fd_sc_hd__nor2_1 _1845_ (.A(\product[13] ),
    .B(\multiplicand[13] ),
    .Y(_0393_));
 sky130_fd_sc_hd__or2_1 _1846_ (.A(\product[13] ),
    .B(\multiplicand[13] ),
    .X(_0394_));
 sky130_fd_sc_hd__and2_1 _1847_ (.A(\product[13] ),
    .B(\multiplicand[13] ),
    .X(_0395_));
 sky130_fd_sc_hd__nor2_1 _1848_ (.A(_0393_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__a22o_2 _1849_ (.A1(\product[12] ),
    .A2(\multiplicand[12] ),
    .B1(\multiplicand[13] ),
    .B2(\product[13] ),
    .X(_0397_));
 sky130_fd_sc_hd__a221o_1 _1850_ (.A1(\product[12] ),
    .A2(\multiplicand[12] ),
    .B1(\multiplicand[13] ),
    .B2(\product[13] ),
    .C1(_0391_),
    .X(_0398_));
 sky130_fd_sc_hd__o22ai_1 _1851_ (.A1(_0386_),
    .A2(_0391_),
    .B1(_0393_),
    .B2(_0395_),
    .Y(_0399_));
 sky130_fd_sc_hd__o2111ai_1 _1852_ (.A1(_0393_),
    .A2(_0398_),
    .B1(_0399_),
    .C1(\multiplier[0] ),
    .D1(_0844_),
    .Y(_0400_));
 sky130_fd_sc_hd__o211a_1 _1853_ (.A1(\product[13] ),
    .A2(net132),
    .B1(_0400_),
    .C1(net142),
    .X(_0172_));
 sky130_fd_sc_hd__nand2_1 _1854_ (.A(\product[14] ),
    .B(\multiplicand[14] ),
    .Y(_0401_));
 sky130_fd_sc_hd__xor2_4 _1855_ (.A(\product[14] ),
    .B(\multiplicand[14] ),
    .X(_0402_));
 sky130_fd_sc_hd__a21o_1 _1856_ (.A1(_0394_),
    .A2(_0398_),
    .B1(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__o221ai_4 _1857_ (.A1(\product[13] ),
    .A2(\multiplicand[13] ),
    .B1(_0397_),
    .B2(_0391_),
    .C1(_0402_),
    .Y(_0404_));
 sky130_fd_sc_hd__a21o_1 _1858_ (.A1(_0403_),
    .A2(_0404_),
    .B1(net131),
    .X(_0405_));
 sky130_fd_sc_hd__o211a_1 _1859_ (.A1(\product[14] ),
    .A2(net132),
    .B1(_0405_),
    .C1(net142),
    .X(_0173_));
 sky130_fd_sc_hd__nor2_1 _1860_ (.A(\product[15] ),
    .B(\multiplicand[15] ),
    .Y(_0406_));
 sky130_fd_sc_hd__and2_1 _1861_ (.A(\product[15] ),
    .B(\multiplicand[15] ),
    .X(_0407_));
 sky130_fd_sc_hd__nor2_2 _1862_ (.A(_0406_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__o2bb2a_1 _1863_ (.A1_N(_0401_),
    .A2_N(_0404_),
    .B1(_0406_),
    .B2(_0407_),
    .X(_0409_));
 sky130_fd_sc_hd__a31o_1 _1864_ (.A1(_0401_),
    .A2(_0404_),
    .A3(_0408_),
    .B1(net131),
    .X(_0410_));
 sky130_fd_sc_hd__o221a_1 _1865_ (.A1(\product[15] ),
    .A2(net132),
    .B1(_0410_),
    .B2(_0409_),
    .C1(net142),
    .X(_0174_));
 sky130_fd_sc_hd__nor2_1 _1866_ (.A(\product[16] ),
    .B(\multiplicand[16] ),
    .Y(_0411_));
 sky130_fd_sc_hd__nand2_1 _1867_ (.A(\product[16] ),
    .B(\multiplicand[16] ),
    .Y(_0412_));
 sky130_fd_sc_hd__and2b_2 _1868_ (.A_N(_0411_),
    .B(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__nand4_4 _1869_ (.A(_0388_),
    .B(_0396_),
    .C(_0402_),
    .D(_0408_),
    .Y(_0414_));
 sky130_fd_sc_hd__nor3_4 _1870_ (.A(_0370_),
    .B(_0380_),
    .C(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__nand4b_2 _1871_ (.A_N(_0414_),
    .B(_0353_),
    .C(_0352_),
    .D(_0384_),
    .Y(_0416_));
 sky130_fd_sc_hd__o21ai_4 _1872_ (.A1(_0349_),
    .A2(_0347_),
    .B1(_0415_),
    .Y(_0417_));
 sky130_fd_sc_hd__o21bai_2 _1873_ (.A1(_0401_),
    .A2(_0406_),
    .B1_N(_0407_),
    .Y(_0418_));
 sky130_fd_sc_hd__a41oi_4 _1874_ (.A1(_0402_),
    .A2(_0408_),
    .A3(_0394_),
    .A4(_0397_),
    .B1(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__o21a_2 _1875_ (.A1(_0414_),
    .A2(_0383_),
    .B1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__o21ai_1 _1876_ (.A1(_0414_),
    .A2(_0383_),
    .B1(_0419_),
    .Y(_0421_));
 sky130_fd_sc_hd__o211a_1 _1877_ (.A1(_0383_),
    .A2(_0414_),
    .B1(_0419_),
    .C1(_0417_),
    .X(_0422_));
 sky130_fd_sc_hd__o21ai_4 _1878_ (.A1(_0416_),
    .A2(net130),
    .B1(_0420_),
    .Y(_0423_));
 sky130_fd_sc_hd__nand2_1 _1879_ (.A(_0423_),
    .B(_0413_),
    .Y(_0424_));
 sky130_fd_sc_hd__a211o_1 _1880_ (.A1(_0351_),
    .A2(_0415_),
    .B1(_0421_),
    .C1(_0413_),
    .X(_0425_));
 sky130_fd_sc_hd__a21oi_1 _1881_ (.A1(_0424_),
    .A2(_0425_),
    .B1(net131),
    .Y(_0426_));
 sky130_fd_sc_hd__a211oi_1 _1882_ (.A1(_0855_),
    .A2(net131),
    .B1(_0426_),
    .C1(net65),
    .Y(_0175_));
 sky130_fd_sc_hd__nor2_1 _1883_ (.A(\product[17] ),
    .B(\multiplicand[17] ),
    .Y(_0427_));
 sky130_fd_sc_hd__and2_1 _1884_ (.A(\product[17] ),
    .B(\multiplicand[17] ),
    .X(_0428_));
 sky130_fd_sc_hd__nand2_1 _1885_ (.A(\product[17] ),
    .B(\multiplicand[17] ),
    .Y(_0429_));
 sky130_fd_sc_hd__nor2_1 _1886_ (.A(_0427_),
    .B(_0428_),
    .Y(_0430_));
 sky130_fd_sc_hd__o2bb2a_1 _1887_ (.A1_N(_0412_),
    .A2_N(_0424_),
    .B1(_0427_),
    .B2(_0428_),
    .X(_0431_));
 sky130_fd_sc_hd__a31o_1 _1888_ (.A1(_0412_),
    .A2(_0424_),
    .A3(_0430_),
    .B1(net131),
    .X(_0432_));
 sky130_fd_sc_hd__o221a_1 _1889_ (.A1(\product[17] ),
    .A2(net132),
    .B1(_0432_),
    .B2(_0431_),
    .C1(net142),
    .X(_0176_));
 sky130_fd_sc_hd__nor2_1 _1890_ (.A(\product[18] ),
    .B(\multiplicand[18] ),
    .Y(_0433_));
 sky130_fd_sc_hd__and2_1 _1891_ (.A(\product[18] ),
    .B(\multiplicand[18] ),
    .X(_0434_));
 sky130_fd_sc_hd__nand2_1 _1892_ (.A(\product[18] ),
    .B(\multiplicand[18] ),
    .Y(_0435_));
 sky130_fd_sc_hd__nor2_1 _1893_ (.A(_0433_),
    .B(_0434_),
    .Y(_0436_));
 sky130_fd_sc_hd__a21oi_1 _1894_ (.A1(_0412_),
    .A2(_0429_),
    .B1(_0427_),
    .Y(_0437_));
 sky130_fd_sc_hd__a31o_1 _1895_ (.A1(_0412_),
    .A2(_0424_),
    .A3(_0429_),
    .B1(_0427_),
    .X(_0438_));
 sky130_fd_sc_hd__nor2_1 _1896_ (.A(_0436_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__a211o_1 _1897_ (.A1(_0436_),
    .A2(_0438_),
    .B1(net131),
    .C1(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__o211a_1 _1898_ (.A1(\product[18] ),
    .A2(net132),
    .B1(_0440_),
    .C1(net142),
    .X(_0177_));
 sky130_fd_sc_hd__nor2_1 _1899_ (.A(\product[19] ),
    .B(\multiplicand[19] ),
    .Y(_0441_));
 sky130_fd_sc_hd__or2_1 _1900_ (.A(\product[19] ),
    .B(\multiplicand[19] ),
    .X(_0442_));
 sky130_fd_sc_hd__and2_1 _1901_ (.A(\product[19] ),
    .B(\multiplicand[19] ),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _1902_ (.A(\product[19] ),
    .B(\multiplicand[19] ),
    .Y(_0444_));
 sky130_fd_sc_hd__nor2_1 _1903_ (.A(_0441_),
    .B(_0443_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_1 _1904_ (.A(_0442_),
    .B(_0444_),
    .Y(_0446_));
 sky130_fd_sc_hd__o21ai_1 _1905_ (.A1(_0433_),
    .A2(_0438_),
    .B1(_0435_),
    .Y(_0447_));
 sky130_fd_sc_hd__o211a_1 _1906_ (.A1(_0433_),
    .A2(_0438_),
    .B1(_0445_),
    .C1(_0435_),
    .X(_0448_));
 sky130_fd_sc_hd__a21o_1 _1907_ (.A1(_0447_),
    .A2(_0446_),
    .B1(net131),
    .X(_0449_));
 sky130_fd_sc_hd__o221a_1 _1908_ (.A1(\product[19] ),
    .A2(net132),
    .B1(_0448_),
    .B2(_0449_),
    .C1(net142),
    .X(_0178_));
 sky130_fd_sc_hd__xor2_2 _1909_ (.A(\product[20] ),
    .B(\multiplicand[20] ),
    .X(_0450_));
 sky130_fd_sc_hd__nand4_2 _1910_ (.A(_0413_),
    .B(_0430_),
    .C(_0436_),
    .D(_0445_),
    .Y(_0451_));
 sky130_fd_sc_hd__nand4_1 _1911_ (.A(_0436_),
    .B(_0437_),
    .C(_0442_),
    .D(_0444_),
    .Y(_0452_));
 sky130_fd_sc_hd__a21o_1 _1912_ (.A1(_0435_),
    .A2(_0444_),
    .B1(_0441_),
    .X(_0453_));
 sky130_fd_sc_hd__o211ai_2 _1913_ (.A1(_0451_),
    .A2(_0422_),
    .B1(_0453_),
    .C1(_0452_),
    .Y(_0454_));
 sky130_fd_sc_hd__nor2_1 _1914_ (.A(_0450_),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_1 _1915_ (.A(_0454_),
    .B(_0450_),
    .Y(_0456_));
 sky130_fd_sc_hd__and2b_1 _1916_ (.A_N(_0455_),
    .B(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__or3b_1 _1917_ (.A(net139),
    .B(_0457_),
    .C_N(\multiplier[0] ),
    .X(_0458_));
 sky130_fd_sc_hd__o211a_1 _1918_ (.A1(\product[20] ),
    .A2(net132),
    .B1(_0458_),
    .C1(net142),
    .X(_0179_));
 sky130_fd_sc_hd__nor2_1 _1919_ (.A(\product[21] ),
    .B(\multiplicand[21] ),
    .Y(_0459_));
 sky130_fd_sc_hd__or2_1 _1920_ (.A(\product[21] ),
    .B(\multiplicand[21] ),
    .X(_0460_));
 sky130_fd_sc_hd__and2_1 _1921_ (.A(\product[21] ),
    .B(\multiplicand[21] ),
    .X(_0461_));
 sky130_fd_sc_hd__nand2_1 _1922_ (.A(\product[21] ),
    .B(\multiplicand[21] ),
    .Y(_0462_));
 sky130_fd_sc_hd__nor2_1 _1923_ (.A(_0459_),
    .B(_0461_),
    .Y(_0463_));
 sky130_fd_sc_hd__a21boi_1 _1924_ (.A1(\product[20] ),
    .A2(\multiplicand[20] ),
    .B1_N(_0456_),
    .Y(_0464_));
 sky130_fd_sc_hd__a21oi_1 _1925_ (.A1(_0460_),
    .A2(_0462_),
    .B1(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__a31o_1 _1926_ (.A1(_0464_),
    .A2(_0462_),
    .A3(_0460_),
    .B1(net131),
    .X(_0466_));
 sky130_fd_sc_hd__o221a_1 _1927_ (.A1(\product[21] ),
    .A2(net132),
    .B1(_0465_),
    .B2(_0466_),
    .C1(net142),
    .X(_0180_));
 sky130_fd_sc_hd__a21oi_1 _1928_ (.A1(\product[20] ),
    .A2(\multiplicand[20] ),
    .B1(_0461_),
    .Y(_0467_));
 sky130_fd_sc_hd__a22o_1 _1929_ (.A1(\product[20] ),
    .A2(\multiplicand[20] ),
    .B1(\multiplicand[21] ),
    .B2(\product[21] ),
    .X(_0468_));
 sky130_fd_sc_hd__a2bb2o_1 _1930_ (.A1_N(\product[21] ),
    .A2_N(\multiplicand[21] ),
    .B1(_0467_),
    .B2(_0456_),
    .X(_0469_));
 sky130_fd_sc_hd__nand2_1 _1931_ (.A(\product[22] ),
    .B(\multiplicand[22] ),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2b_1 _1932_ (.A_N(\product[22] ),
    .B(\multiplicand[22] ),
    .Y(_0471_));
 sky130_fd_sc_hd__nand2b_1 _1933_ (.A_N(\multiplicand[22] ),
    .B(\product[22] ),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_2 _1934_ (.A(_0471_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__a221o_1 _1935_ (.A1(_0471_),
    .A2(_0472_),
    .B1(_0456_),
    .B2(_0467_),
    .C1(_0459_),
    .X(_0474_));
 sky130_fd_sc_hd__xnor2_1 _1936_ (.A(_0469_),
    .B(_0473_),
    .Y(_0475_));
 sky130_fd_sc_hd__a21o_1 _1937_ (.A1(_0844_),
    .A2(\multiplier[0] ),
    .B1(\product[22] ),
    .X(_0476_));
 sky130_fd_sc_hd__o211a_1 _1938_ (.A1(net131),
    .A2(_0475_),
    .B1(_0476_),
    .C1(net142),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_1 _1939_ (.A(\product[23] ),
    .B(\multiplicand[23] ),
    .Y(_0477_));
 sky130_fd_sc_hd__nor2_1 _1940_ (.A(\product[23] ),
    .B(\multiplicand[23] ),
    .Y(_0478_));
 sky130_fd_sc_hd__nand2b_1 _1941_ (.A_N(\product[23] ),
    .B(\multiplicand[23] ),
    .Y(_0479_));
 sky130_fd_sc_hd__nand2b_1 _1942_ (.A_N(\multiplicand[23] ),
    .B(\product[23] ),
    .Y(_0480_));
 sky130_fd_sc_hd__nand2_2 _1943_ (.A(_0479_),
    .B(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__a21oi_1 _1944_ (.A1(_0470_),
    .A2(_0474_),
    .B1(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__a31o_1 _1945_ (.A1(_0470_),
    .A2(_0474_),
    .A3(_0481_),
    .B1(net131),
    .X(_0483_));
 sky130_fd_sc_hd__o221a_1 _1946_ (.A1(\product[23] ),
    .A2(net132),
    .B1(_0482_),
    .B2(_0483_),
    .C1(net142),
    .X(_0182_));
 sky130_fd_sc_hd__nor2_1 _1947_ (.A(\product[24] ),
    .B(\multiplicand[24] ),
    .Y(_0484_));
 sky130_fd_sc_hd__and2_1 _1948_ (.A(\product[24] ),
    .B(\multiplicand[24] ),
    .X(_0485_));
 sky130_fd_sc_hd__nand2_1 _1949_ (.A(\product[24] ),
    .B(\multiplicand[24] ),
    .Y(_0486_));
 sky130_fd_sc_hd__nand4_2 _1950_ (.A(_0450_),
    .B(_0463_),
    .C(_0473_),
    .D(_0481_),
    .Y(_0487_));
 sky130_fd_sc_hd__nor2_2 _1951_ (.A(_0451_),
    .B(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__a21oi_1 _1952_ (.A1(_0452_),
    .A2(_0453_),
    .B1(_0487_),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_1 _1953_ (.A1(_0470_),
    .A2(_0478_),
    .B1(_0477_),
    .Y(_0490_));
 sky130_fd_sc_hd__a41o_1 _1954_ (.A1(_0473_),
    .A2(_0481_),
    .A3(_0460_),
    .A4(_0468_),
    .B1(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__or2_1 _1955_ (.A(_0491_),
    .B(_0489_),
    .X(_0492_));
 sky130_fd_sc_hd__a21oi_4 _1956_ (.A1(_0423_),
    .A2(_0488_),
    .B1(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__o21ai_1 _1957_ (.A1(_0484_),
    .A2(_0485_),
    .B1(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__or3_1 _1958_ (.A(_0484_),
    .B(_0485_),
    .C(_0493_),
    .X(_0495_));
 sky130_fd_sc_hd__a21o_1 _1959_ (.A1(_0494_),
    .A2(_0495_),
    .B1(net131),
    .X(_0496_));
 sky130_fd_sc_hd__o211a_1 _1960_ (.A1(\product[24] ),
    .A2(net132),
    .B1(_0496_),
    .C1(net142),
    .X(_0183_));
 sky130_fd_sc_hd__nor2_1 _1961_ (.A(\product[25] ),
    .B(\multiplicand[25] ),
    .Y(_0497_));
 sky130_fd_sc_hd__or2_1 _1962_ (.A(\product[25] ),
    .B(\multiplicand[25] ),
    .X(_0498_));
 sky130_fd_sc_hd__nand2_1 _1963_ (.A(\product[25] ),
    .B(\multiplicand[25] ),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _1964_ (.A(_0498_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__o21ai_1 _1965_ (.A1(_0484_),
    .A2(_0493_),
    .B1(_0486_),
    .Y(_0501_));
 sky130_fd_sc_hd__o2111a_1 _1966_ (.A1(_0484_),
    .A2(_0493_),
    .B1(_0498_),
    .C1(_0499_),
    .D1(_0486_),
    .X(_0502_));
 sky130_fd_sc_hd__a21o_1 _1967_ (.A1(_0500_),
    .A2(_0501_),
    .B1(net131),
    .X(_0503_));
 sky130_fd_sc_hd__o221a_1 _1968_ (.A1(\product[25] ),
    .A2(net132),
    .B1(_0502_),
    .B2(_0503_),
    .C1(net142),
    .X(_0184_));
 sky130_fd_sc_hd__or2_1 _1969_ (.A(\product[26] ),
    .B(\multiplicand[26] ),
    .X(_0504_));
 sky130_fd_sc_hd__nand2_2 _1970_ (.A(\product[26] ),
    .B(\multiplicand[26] ),
    .Y(_0505_));
 sky130_fd_sc_hd__nand2_1 _1971_ (.A(_0504_),
    .B(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__o21ai_1 _1972_ (.A1(_0486_),
    .A2(_0497_),
    .B1(_0499_),
    .Y(_0507_));
 sky130_fd_sc_hd__nand4b_2 _1973_ (.A_N(_0484_),
    .B(_0486_),
    .C(_0498_),
    .D(_0499_),
    .Y(_0508_));
 sky130_fd_sc_hd__o21bai_2 _1974_ (.A1(_0508_),
    .A2(_0493_),
    .B1_N(_0507_),
    .Y(_0509_));
 sky130_fd_sc_hd__a21oi_1 _1975_ (.A1(_0506_),
    .A2(_0509_),
    .B1(net131),
    .Y(_0510_));
 sky130_fd_sc_hd__o21ai_1 _1976_ (.A1(_0506_),
    .A2(_0509_),
    .B1(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__o211a_1 _1977_ (.A1(\product[26] ),
    .A2(net132),
    .B1(_0511_),
    .C1(net142),
    .X(_0185_));
 sky130_fd_sc_hd__nor2_1 _1978_ (.A(\product[27] ),
    .B(\multiplicand[27] ),
    .Y(_0512_));
 sky130_fd_sc_hd__and2_1 _1979_ (.A(\product[27] ),
    .B(\multiplicand[27] ),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _1980_ (.A(\product[27] ),
    .B(\multiplicand[27] ),
    .Y(_0514_));
 sky130_fd_sc_hd__nor2_1 _1981_ (.A(_0512_),
    .B(_0513_),
    .Y(_0515_));
 sky130_fd_sc_hd__o21ai_1 _1982_ (.A1(\product[26] ),
    .A2(\multiplicand[26] ),
    .B1(_0509_),
    .Y(_0516_));
 sky130_fd_sc_hd__a21oi_1 _1983_ (.A1(_0505_),
    .A2(_0516_),
    .B1(_0515_),
    .Y(_0517_));
 sky130_fd_sc_hd__a31o_1 _1984_ (.A1(_0505_),
    .A2(_0516_),
    .A3(_0515_),
    .B1(net131),
    .X(_0518_));
 sky130_fd_sc_hd__o221a_1 _1985_ (.A1(\product[27] ),
    .A2(net132),
    .B1(_0517_),
    .B2(_0518_),
    .C1(net142),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _1986_ (.A(_0515_),
    .B(_0505_),
    .C(_0504_),
    .X(_0519_));
 sky130_fd_sc_hd__nand3_1 _1987_ (.A(_0515_),
    .B(_0505_),
    .C(_0504_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2_1 _1988_ (.A(_0509_),
    .B(_0519_),
    .Y(_0521_));
 sky130_fd_sc_hd__a21o_1 _1989_ (.A1(_0505_),
    .A2(_0514_),
    .B1(_0512_),
    .X(_0522_));
 sky130_fd_sc_hd__a21oi_1 _1990_ (.A1(_0505_),
    .A2(_0514_),
    .B1(_0512_),
    .Y(_0523_));
 sky130_fd_sc_hd__xor2_1 _1991_ (.A(\product[28] ),
    .B(\multiplicand[28] ),
    .X(_0524_));
 sky130_fd_sc_hd__xnor2_2 _1992_ (.A(\product[28] ),
    .B(\multiplicand[28] ),
    .Y(_0525_));
 sky130_fd_sc_hd__and3_1 _1993_ (.A(_0521_),
    .B(_0522_),
    .C(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__a21oi_4 _1994_ (.A1(_0521_),
    .A2(_0522_),
    .B1(_0525_),
    .Y(_0527_));
 sky130_fd_sc_hd__o21ai_1 _1995_ (.A1(_0526_),
    .A2(_0527_),
    .B1(net132),
    .Y(_0528_));
 sky130_fd_sc_hd__o211a_1 _1996_ (.A1(\product[28] ),
    .A2(net132),
    .B1(_0528_),
    .C1(net142),
    .X(_0187_));
 sky130_fd_sc_hd__nor2_1 _1997_ (.A(\product[29] ),
    .B(\multiplicand[29] ),
    .Y(_0529_));
 sky130_fd_sc_hd__and2_1 _1998_ (.A(\product[29] ),
    .B(\multiplicand[29] ),
    .X(_0530_));
 sky130_fd_sc_hd__nor2_1 _1999_ (.A(_0529_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__a21oi_1 _2000_ (.A1(\product[28] ),
    .A2(\multiplicand[28] ),
    .B1(_0527_),
    .Y(_0532_));
 sky130_fd_sc_hd__a22o_2 _2001_ (.A1(\product[28] ),
    .A2(\multiplicand[28] ),
    .B1(\multiplicand[29] ),
    .B2(\product[29] ),
    .X(_0533_));
 sky130_fd_sc_hd__or2_1 _2002_ (.A(_0531_),
    .B(_0532_),
    .X(_0534_));
 sky130_fd_sc_hd__o311a_1 _2003_ (.A1(_0533_),
    .A2(_0529_),
    .A3(_0527_),
    .B1(_0844_),
    .C1(\multiplier[0] ),
    .X(_0535_));
 sky130_fd_sc_hd__a21oi_1 _2004_ (.A1(_0844_),
    .A2(\multiplier[0] ),
    .B1(\product[29] ),
    .Y(_0536_));
 sky130_fd_sc_hd__a211oi_1 _2005_ (.A1(_0534_),
    .A2(_0535_),
    .B1(_0536_),
    .C1(net65),
    .Y(_0188_));
 sky130_fd_sc_hd__nor2_1 _2006_ (.A(\product[30] ),
    .B(\multiplicand[30] ),
    .Y(_0537_));
 sky130_fd_sc_hd__and2_1 _2007_ (.A(\product[30] ),
    .B(\multiplicand[30] ),
    .X(_0538_));
 sky130_fd_sc_hd__nor2_1 _2008_ (.A(_0537_),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__o22ai_1 _2009_ (.A1(\product[29] ),
    .A2(\multiplicand[29] ),
    .B1(_0533_),
    .B2(_0527_),
    .Y(_0540_));
 sky130_fd_sc_hd__o21ai_1 _2010_ (.A1(_0537_),
    .A2(_0538_),
    .B1(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__o221a_1 _2011_ (.A1(\product[29] ),
    .A2(\multiplicand[29] ),
    .B1(_0533_),
    .B2(_0527_),
    .C1(_0539_),
    .X(_0542_));
 sky130_fd_sc_hd__o221ai_2 _2012_ (.A1(\product[29] ),
    .A2(\multiplicand[29] ),
    .B1(_0533_),
    .B2(_0527_),
    .C1(_0539_),
    .Y(_0543_));
 sky130_fd_sc_hd__a21o_1 _2013_ (.A1(_0541_),
    .A2(_0543_),
    .B1(net131),
    .X(_0544_));
 sky130_fd_sc_hd__o211a_1 _2014_ (.A1(\product[30] ),
    .A2(net132),
    .B1(_0544_),
    .C1(net142),
    .X(_0189_));
 sky130_fd_sc_hd__nor2_1 _2015_ (.A(\product[31] ),
    .B(\multiplicand[31] ),
    .Y(_0545_));
 sky130_fd_sc_hd__and2_1 _2016_ (.A(\product[31] ),
    .B(\multiplicand[31] ),
    .X(_0546_));
 sky130_fd_sc_hd__nor2_1 _2017_ (.A(_0545_),
    .B(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__o22ai_1 _2018_ (.A1(_0538_),
    .A2(_0542_),
    .B1(_0545_),
    .B2(_0546_),
    .Y(_0548_));
 sky130_fd_sc_hd__nand3b_1 _2019_ (.A_N(_0538_),
    .B(_0543_),
    .C(_0547_),
    .Y(_0549_));
 sky130_fd_sc_hd__o21ai_1 _2020_ (.A1(\product[31] ),
    .A2(net132),
    .B1(net142),
    .Y(_0550_));
 sky130_fd_sc_hd__a31oi_1 _2021_ (.A1(_0548_),
    .A2(_0549_),
    .A3(net132),
    .B1(_0550_),
    .Y(_0190_));
 sky130_fd_sc_hd__or2_1 _2022_ (.A(\product[32] ),
    .B(\multiplicand[32] ),
    .X(_0551_));
 sky130_fd_sc_hd__nand2_1 _2023_ (.A(\product[32] ),
    .B(\multiplicand[32] ),
    .Y(_0552_));
 sky130_fd_sc_hd__nand2_1 _2024_ (.A(_0551_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__nand2_1 _2025_ (.A(_0524_),
    .B(_0531_),
    .Y(_0554_));
 sky130_fd_sc_hd__nand4_1 _2026_ (.A(_0524_),
    .B(_0531_),
    .C(_0539_),
    .D(_0547_),
    .Y(_0555_));
 sky130_fd_sc_hd__nor3_2 _2027_ (.A(_0508_),
    .B(_0520_),
    .C(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__and2_4 _2028_ (.A(_0488_),
    .B(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__nand2_2 _2029_ (.A(_0488_),
    .B(_0556_),
    .Y(_0558_));
 sky130_fd_sc_hd__a21oi_4 _2030_ (.A1(_0417_),
    .A2(_0420_),
    .B1(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__a41oi_2 _2031_ (.A1(_0515_),
    .A2(_0507_),
    .A3(_0505_),
    .A4(_0504_),
    .B1(_0523_),
    .Y(_0560_));
 sky130_fd_sc_hd__o21ai_1 _2032_ (.A1(\product[29] ),
    .A2(\multiplicand[29] ),
    .B1(_0533_),
    .Y(_0561_));
 sky130_fd_sc_hd__o21ai_1 _2033_ (.A1(_0554_),
    .A2(_0560_),
    .B1(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand3_1 _2034_ (.A(_0562_),
    .B(_0547_),
    .C(_0539_),
    .Y(_0563_));
 sky130_fd_sc_hd__o21ai_2 _2035_ (.A1(_0491_),
    .A2(_0489_),
    .B1(_0556_),
    .Y(_0564_));
 sky130_fd_sc_hd__o21bai_2 _2036_ (.A1(_0538_),
    .A2(_0546_),
    .B1_N(_0545_),
    .Y(_0565_));
 sky130_fd_sc_hd__nand3_4 _2037_ (.A(_0563_),
    .B(_0564_),
    .C(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__a21oi_4 _2038_ (.A1(_0423_),
    .A2(_0557_),
    .B1(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__o211a_1 _2039_ (.A1(_0566_),
    .A2(_0559_),
    .B1(_0552_),
    .C1(_0551_),
    .X(_0568_));
 sky130_fd_sc_hd__a221oi_1 _2040_ (.A1(_0551_),
    .A2(_0552_),
    .B1(_0423_),
    .B2(_0557_),
    .C1(_0566_),
    .Y(_0569_));
 sky130_fd_sc_hd__o21ai_1 _2041_ (.A1(_0568_),
    .A2(_0569_),
    .B1(net132),
    .Y(_0570_));
 sky130_fd_sc_hd__o211a_1 _2042_ (.A1(\product[32] ),
    .A2(net132),
    .B1(_0570_),
    .C1(_0859_),
    .X(_0191_));
 sky130_fd_sc_hd__o21ai_1 _2043_ (.A1(_0553_),
    .A2(_0567_),
    .B1(_0552_),
    .Y(_0571_));
 sky130_fd_sc_hd__nor2_1 _2044_ (.A(\product[33] ),
    .B(\multiplicand[33] ),
    .Y(_0572_));
 sky130_fd_sc_hd__and2_1 _2045_ (.A(\product[33] ),
    .B(\multiplicand[33] ),
    .X(_0573_));
 sky130_fd_sc_hd__o21a_1 _2046_ (.A1(_0572_),
    .A2(_0573_),
    .B1(_0571_),
    .X(_0574_));
 sky130_fd_sc_hd__o31ai_1 _2047_ (.A1(_0572_),
    .A2(_0573_),
    .A3(_0571_),
    .B1(net132),
    .Y(_0575_));
 sky130_fd_sc_hd__o221a_1 _2048_ (.A1(\product[33] ),
    .A2(net132),
    .B1(_0574_),
    .B2(_0575_),
    .C1(_0859_),
    .X(_0192_));
 sky130_fd_sc_hd__a22o_1 _2049_ (.A1(\product[32] ),
    .A2(\multiplicand[32] ),
    .B1(\multiplicand[33] ),
    .B2(\product[33] ),
    .X(_0576_));
 sky130_fd_sc_hd__o21ai_1 _2050_ (.A1(\product[33] ),
    .A2(\multiplicand[33] ),
    .B1(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__o21a_1 _2051_ (.A1(\product[33] ),
    .A2(\multiplicand[33] ),
    .B1(_0576_),
    .X(_0578_));
 sky130_fd_sc_hd__o31a_1 _2052_ (.A1(_0572_),
    .A2(_0553_),
    .A3(_0567_),
    .B1(_0577_),
    .X(_0579_));
 sky130_fd_sc_hd__and2_1 _2053_ (.A(\product[34] ),
    .B(\multiplicand[34] ),
    .X(_0580_));
 sky130_fd_sc_hd__nor2_1 _2054_ (.A(\product[34] ),
    .B(\multiplicand[34] ),
    .Y(_0581_));
 sky130_fd_sc_hd__nor2_1 _2055_ (.A(_0580_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__xnor2_1 _2056_ (.A(_0579_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__a21o_1 _2057_ (.A1(_0844_),
    .A2(\multiplier[0] ),
    .B1(\product[34] ),
    .X(_0584_));
 sky130_fd_sc_hd__o211a_1 _2058_ (.A1(_0288_),
    .A2(_0583_),
    .B1(_0584_),
    .C1(_0859_),
    .X(_0193_));
 sky130_fd_sc_hd__nor2_1 _2059_ (.A(\product[35] ),
    .B(\multiplicand[35] ),
    .Y(_0585_));
 sky130_fd_sc_hd__and2_1 _2060_ (.A(\product[35] ),
    .B(\multiplicand[35] ),
    .X(_0586_));
 sky130_fd_sc_hd__nor2_1 _2061_ (.A(_0585_),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__o21bai_1 _2062_ (.A1(_0579_),
    .A2(_0581_),
    .B1_N(_0580_),
    .Y(_0588_));
 sky130_fd_sc_hd__o21a_1 _2063_ (.A1(_0585_),
    .A2(_0586_),
    .B1(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__o31ai_1 _2064_ (.A1(_0585_),
    .A2(_0586_),
    .A3(_0588_),
    .B1(net132),
    .Y(_0590_));
 sky130_fd_sc_hd__o221a_1 _2065_ (.A1(\product[35] ),
    .A2(net132),
    .B1(_0589_),
    .B2(_0590_),
    .C1(_0859_),
    .X(_0194_));
 sky130_fd_sc_hd__nor2_1 _2066_ (.A(\product[36] ),
    .B(\multiplicand[36] ),
    .Y(_0591_));
 sky130_fd_sc_hd__and2_1 _2067_ (.A(\product[36] ),
    .B(\multiplicand[36] ),
    .X(_0592_));
 sky130_fd_sc_hd__nor2_2 _2068_ (.A(_0591_),
    .B(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__o21ba_1 _2069_ (.A1(_0580_),
    .A2(_0586_),
    .B1_N(_0585_),
    .X(_0594_));
 sky130_fd_sc_hd__a31oi_2 _2070_ (.A1(_0578_),
    .A2(_0582_),
    .A3(_0587_),
    .B1(_0594_),
    .Y(_0595_));
 sky130_fd_sc_hd__nor3_1 _2071_ (.A(_0572_),
    .B(_0573_),
    .C(_0553_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand3_2 _2072_ (.A(_0582_),
    .B(_0587_),
    .C(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__o21ai_2 _2073_ (.A1(_0597_),
    .A2(_0567_),
    .B1(_0595_),
    .Y(_0598_));
 sky130_fd_sc_hd__xor2_1 _2074_ (.A(_0593_),
    .B(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__or3b_1 _2075_ (.A(net141),
    .B(_0599_),
    .C_N(\multiplier[0] ),
    .X(_0600_));
 sky130_fd_sc_hd__o211a_1 _2076_ (.A1(\product[36] ),
    .A2(net132),
    .B1(_0600_),
    .C1(_0859_),
    .X(_0195_));
 sky130_fd_sc_hd__a21oi_1 _2077_ (.A1(_0598_),
    .A2(_0593_),
    .B1(_0592_),
    .Y(_0601_));
 sky130_fd_sc_hd__nor2_1 _2078_ (.A(\product[37] ),
    .B(\multiplicand[37] ),
    .Y(_0602_));
 sky130_fd_sc_hd__and2_1 _2079_ (.A(\product[37] ),
    .B(\multiplicand[37] ),
    .X(_0603_));
 sky130_fd_sc_hd__nor2_1 _2080_ (.A(_0602_),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__a22o_1 _2081_ (.A1(\product[36] ),
    .A2(\multiplicand[36] ),
    .B1(\multiplicand[37] ),
    .B2(\product[37] ),
    .X(_0605_));
 sky130_fd_sc_hd__a21oi_2 _2082_ (.A1(_0598_),
    .A2(_0593_),
    .B1(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__o21a_1 _2083_ (.A1(\product[37] ),
    .A2(\multiplicand[37] ),
    .B1(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__o21ai_1 _2084_ (.A1(_0601_),
    .A2(_0604_),
    .B1(net132),
    .Y(_0608_));
 sky130_fd_sc_hd__o221a_1 _2085_ (.A1(\product[37] ),
    .A2(net132),
    .B1(_0607_),
    .B2(_0608_),
    .C1(_0859_),
    .X(_0196_));
 sky130_fd_sc_hd__nor2_1 _2086_ (.A(\product[38] ),
    .B(\multiplicand[38] ),
    .Y(_0609_));
 sky130_fd_sc_hd__nand2_1 _2087_ (.A(\product[38] ),
    .B(\multiplicand[38] ),
    .Y(_0610_));
 sky130_fd_sc_hd__and2b_1 _2088_ (.A_N(_0609_),
    .B(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__o21ba_1 _2089_ (.A1(_0602_),
    .A2(_0606_),
    .B1_N(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__nor4b_1 _2090_ (.A(_0602_),
    .B(_0606_),
    .C(_0609_),
    .D_N(_0610_),
    .Y(_0613_));
 sky130_fd_sc_hd__o21ai_1 _2091_ (.A1(_0612_),
    .A2(_0613_),
    .B1(net132),
    .Y(_0614_));
 sky130_fd_sc_hd__o211a_1 _2092_ (.A1(\product[38] ),
    .A2(net132),
    .B1(_0614_),
    .C1(_0859_),
    .X(_0197_));
 sky130_fd_sc_hd__o31ai_1 _2093_ (.A1(_0602_),
    .A2(_0606_),
    .A3(_0609_),
    .B1(_0610_),
    .Y(_0615_));
 sky130_fd_sc_hd__xor2_1 _2094_ (.A(\product[39] ),
    .B(\multiplicand[39] ),
    .X(_0616_));
 sky130_fd_sc_hd__xnor2_1 _2095_ (.A(\product[39] ),
    .B(\multiplicand[39] ),
    .Y(_0617_));
 sky130_fd_sc_hd__a21oi_1 _2096_ (.A1(_0615_),
    .A2(_0617_),
    .B1(_0288_),
    .Y(_0618_));
 sky130_fd_sc_hd__o21ai_1 _2097_ (.A1(_0615_),
    .A2(_0617_),
    .B1(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__o211a_1 _2098_ (.A1(\product[39] ),
    .A2(net132),
    .B1(_0619_),
    .C1(_0859_),
    .X(_0198_));
 sky130_fd_sc_hd__or2_1 _2099_ (.A(\product[40] ),
    .B(\multiplicand[40] ),
    .X(_0620_));
 sky130_fd_sc_hd__nand2_1 _2100_ (.A(\product[40] ),
    .B(\multiplicand[40] ),
    .Y(_0621_));
 sky130_fd_sc_hd__and2_1 _2101_ (.A(_0620_),
    .B(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__nand4_2 _2102_ (.A(_0593_),
    .B(_0604_),
    .C(_0611_),
    .D(_0616_),
    .Y(_0623_));
 sky130_fd_sc_hd__o2111ai_1 _2103_ (.A1(\product[37] ),
    .A2(\multiplicand[37] ),
    .B1(_0605_),
    .C1(_0611_),
    .D1(_0616_),
    .Y(_0624_));
 sky130_fd_sc_hd__o211a_1 _2104_ (.A1(\product[39] ),
    .A2(\multiplicand[39] ),
    .B1(\multiplicand[38] ),
    .C1(\product[38] ),
    .X(_0625_));
 sky130_fd_sc_hd__a21oi_1 _2105_ (.A1(\product[39] ),
    .A2(\multiplicand[39] ),
    .B1(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__o211a_1 _2106_ (.A1(_0623_),
    .A2(_0595_),
    .B1(_0626_),
    .C1(_0624_),
    .X(_0627_));
 sky130_fd_sc_hd__nor2_1 _2107_ (.A(_0597_),
    .B(_0623_),
    .Y(_0628_));
 sky130_fd_sc_hd__or2_1 _2108_ (.A(_0597_),
    .B(_0623_),
    .X(_0629_));
 sky130_fd_sc_hd__o21ai_1 _2109_ (.A1(_0566_),
    .A2(_0559_),
    .B1(_0628_),
    .Y(_0630_));
 sky130_fd_sc_hd__o21ai_1 _2110_ (.A1(_0629_),
    .A2(_0567_),
    .B1(_0627_),
    .Y(_0631_));
 sky130_fd_sc_hd__nand2_1 _2111_ (.A(_0631_),
    .B(_0622_),
    .Y(_0632_));
 sky130_fd_sc_hd__xor2_1 _2112_ (.A(_0622_),
    .B(_0631_),
    .X(_0633_));
 sky130_fd_sc_hd__or3b_1 _2113_ (.A(net140),
    .B(_0633_),
    .C_N(\multiplier[0] ),
    .X(_0634_));
 sky130_fd_sc_hd__o211a_1 _2114_ (.A1(\product[40] ),
    .A2(net133),
    .B1(_0634_),
    .C1(_0859_),
    .X(_0199_));
 sky130_fd_sc_hd__nor2_1 _2115_ (.A(\product[41] ),
    .B(\multiplicand[41] ),
    .Y(_0635_));
 sky130_fd_sc_hd__or2_1 _2116_ (.A(\product[41] ),
    .B(\multiplicand[41] ),
    .X(_0636_));
 sky130_fd_sc_hd__and2_1 _2117_ (.A(\product[41] ),
    .B(\multiplicand[41] ),
    .X(_0637_));
 sky130_fd_sc_hd__nor2_1 _2118_ (.A(_0635_),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__o2bb2a_1 _2119_ (.A1_N(_0621_),
    .A2_N(_0632_),
    .B1(_0635_),
    .B2(_0637_),
    .X(_0639_));
 sky130_fd_sc_hd__a31o_1 _2120_ (.A1(_0621_),
    .A2(_0632_),
    .A3(_0638_),
    .B1(_0288_),
    .X(_0640_));
 sky130_fd_sc_hd__o221a_1 _2121_ (.A1(\product[41] ),
    .A2(net133),
    .B1(_0639_),
    .B2(_0640_),
    .C1(_0859_),
    .X(_0200_));
 sky130_fd_sc_hd__or2_1 _2122_ (.A(\product[42] ),
    .B(\multiplicand[42] ),
    .X(_0641_));
 sky130_fd_sc_hd__nand2_2 _2123_ (.A(\product[42] ),
    .B(\multiplicand[42] ),
    .Y(_0642_));
 sky130_fd_sc_hd__and2_1 _2124_ (.A(_0641_),
    .B(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__a21oi_1 _2125_ (.A1(\product[40] ),
    .A2(\multiplicand[40] ),
    .B1(_0637_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_1 _2126_ (.A(_0632_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__a22o_1 _2127_ (.A1(_0641_),
    .A2(_0642_),
    .B1(_0645_),
    .B2(_0636_),
    .X(_0646_));
 sky130_fd_sc_hd__o2111ai_4 _2128_ (.A1(\product[41] ),
    .A2(\multiplicand[41] ),
    .B1(_0641_),
    .C1(_0642_),
    .D1(_0645_),
    .Y(_0647_));
 sky130_fd_sc_hd__a21o_1 _2129_ (.A1(_0646_),
    .A2(_0647_),
    .B1(_0288_),
    .X(_0648_));
 sky130_fd_sc_hd__o211a_1 _2130_ (.A1(\product[42] ),
    .A2(net133),
    .B1(_0648_),
    .C1(_0859_),
    .X(_0201_));
 sky130_fd_sc_hd__nor2_1 _2131_ (.A(\product[43] ),
    .B(\multiplicand[43] ),
    .Y(_0649_));
 sky130_fd_sc_hd__and2_1 _2132_ (.A(\product[43] ),
    .B(\multiplicand[43] ),
    .X(_0650_));
 sky130_fd_sc_hd__nor2_1 _2133_ (.A(_0649_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__o2bb2a_1 _2134_ (.A1_N(_0642_),
    .A2_N(_0647_),
    .B1(_0649_),
    .B2(_0650_),
    .X(_0652_));
 sky130_fd_sc_hd__a31o_1 _2135_ (.A1(_0642_),
    .A2(_0647_),
    .A3(_0651_),
    .B1(_0288_),
    .X(_0653_));
 sky130_fd_sc_hd__o221a_1 _2136_ (.A1(\product[43] ),
    .A2(net133),
    .B1(_0653_),
    .B2(_0652_),
    .C1(_0859_),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _2137_ (.A(\product[44] ),
    .B(\multiplicand[44] ),
    .X(_0654_));
 sky130_fd_sc_hd__nand2_1 _2138_ (.A(\product[44] ),
    .B(\multiplicand[44] ),
    .Y(_0655_));
 sky130_fd_sc_hd__nor2_1 _2139_ (.A(\product[44] ),
    .B(\multiplicand[44] ),
    .Y(_0656_));
 sky130_fd_sc_hd__nor2_1 _2140_ (.A(_0654_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__nand2_1 _2141_ (.A(_0643_),
    .B(_0651_),
    .Y(_0658_));
 sky130_fd_sc_hd__nand4_2 _2142_ (.A(_0622_),
    .B(_0638_),
    .C(_0643_),
    .D(_0651_),
    .Y(_0659_));
 sky130_fd_sc_hd__a21oi_1 _2143_ (.A1(_0630_),
    .A2(_0627_),
    .B1(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__a21oi_1 _2144_ (.A1(\product[42] ),
    .A2(\multiplicand[42] ),
    .B1(_0650_),
    .Y(_0661_));
 sky130_fd_sc_hd__o32a_1 _2145_ (.A1(_0635_),
    .A2(_0644_),
    .A3(_0658_),
    .B1(_0661_),
    .B2(_0649_),
    .X(_0662_));
 sky130_fd_sc_hd__inv_2 _2146_ (.A(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__o21ai_1 _2147_ (.A1(_0654_),
    .A2(_0656_),
    .B1(_0662_),
    .Y(_0664_));
 sky130_fd_sc_hd__o21ai_2 _2148_ (.A1(_0663_),
    .A2(_0660_),
    .B1(_0657_),
    .Y(_0665_));
 sky130_fd_sc_hd__o21a_1 _2149_ (.A1(_0660_),
    .A2(_0664_),
    .B1(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__a21o_1 _2150_ (.A1(_0844_),
    .A2(\multiplier[0] ),
    .B1(\product[44] ),
    .X(_0667_));
 sky130_fd_sc_hd__o211a_1 _2151_ (.A1(_0288_),
    .A2(_0666_),
    .B1(_0667_),
    .C1(_0859_),
    .X(_0203_));
 sky130_fd_sc_hd__or2_1 _2152_ (.A(\product[45] ),
    .B(\multiplicand[45] ),
    .X(_0668_));
 sky130_fd_sc_hd__nand2_1 _2153_ (.A(\product[45] ),
    .B(\multiplicand[45] ),
    .Y(_0669_));
 sky130_fd_sc_hd__and2_1 _2154_ (.A(_0668_),
    .B(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__a21oi_1 _2155_ (.A1(_0655_),
    .A2(_0665_),
    .B1(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__a31o_1 _2156_ (.A1(_0655_),
    .A2(_0665_),
    .A3(_0670_),
    .B1(_0288_),
    .X(_0672_));
 sky130_fd_sc_hd__o221a_1 _2157_ (.A1(\product[45] ),
    .A2(net133),
    .B1(_0671_),
    .B2(_0672_),
    .C1(_0859_),
    .X(_0204_));
 sky130_fd_sc_hd__and2_1 _2158_ (.A(\product[46] ),
    .B(\multiplicand[46] ),
    .X(_0673_));
 sky130_fd_sc_hd__nor2_1 _2159_ (.A(\product[46] ),
    .B(\multiplicand[46] ),
    .Y(_0674_));
 sky130_fd_sc_hd__nor2_1 _2160_ (.A(_0673_),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__a21oi_1 _2161_ (.A1(\product[45] ),
    .A2(\multiplicand[45] ),
    .B1(_0654_),
    .Y(_0676_));
 sky130_fd_sc_hd__a22o_1 _2162_ (.A1(\product[44] ),
    .A2(\multiplicand[44] ),
    .B1(\multiplicand[45] ),
    .B2(\product[45] ),
    .X(_0677_));
 sky130_fd_sc_hd__nand2_1 _2163_ (.A(_0665_),
    .B(_0676_),
    .Y(_0678_));
 sky130_fd_sc_hd__a21oi_1 _2164_ (.A1(_0668_),
    .A2(_0678_),
    .B1(_0675_),
    .Y(_0679_));
 sky130_fd_sc_hd__o21ai_1 _2165_ (.A1(\product[45] ),
    .A2(\multiplicand[45] ),
    .B1(_0675_),
    .Y(_0680_));
 sky130_fd_sc_hd__a21oi_1 _2166_ (.A1(_0665_),
    .A2(_0676_),
    .B1(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__o21ai_1 _2167_ (.A1(_0679_),
    .A2(_0681_),
    .B1(net133),
    .Y(_0682_));
 sky130_fd_sc_hd__o211a_1 _2168_ (.A1(\product[46] ),
    .A2(net133),
    .B1(_0682_),
    .C1(_0859_),
    .X(_0205_));
 sky130_fd_sc_hd__a21oi_1 _2169_ (.A1(\product[46] ),
    .A2(\multiplicand[46] ),
    .B1(_0681_),
    .Y(_0683_));
 sky130_fd_sc_hd__xor2_2 _2170_ (.A(\product[47] ),
    .B(\multiplicand[47] ),
    .X(_0684_));
 sky130_fd_sc_hd__o21bai_1 _2171_ (.A1(_0673_),
    .A2(_0681_),
    .B1_N(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__nand2_1 _2172_ (.A(_0683_),
    .B(_0684_),
    .Y(_0686_));
 sky130_fd_sc_hd__a21oi_1 _2173_ (.A1(_0844_),
    .A2(\multiplier[0] ),
    .B1(\product[47] ),
    .Y(_0687_));
 sky130_fd_sc_hd__a311oi_1 _2174_ (.A1(_0686_),
    .A2(net133),
    .A3(_0685_),
    .B1(_0687_),
    .C1(net65),
    .Y(_0206_));
 sky130_fd_sc_hd__nor2_1 _2175_ (.A(\product[48] ),
    .B(\multiplicand[48] ),
    .Y(_0688_));
 sky130_fd_sc_hd__and2_1 _2176_ (.A(\product[48] ),
    .B(\multiplicand[48] ),
    .X(_0689_));
 sky130_fd_sc_hd__nand2_1 _2177_ (.A(\product[48] ),
    .B(\multiplicand[48] ),
    .Y(_0690_));
 sky130_fd_sc_hd__nor2_1 _2178_ (.A(_0688_),
    .B(_0689_),
    .Y(_0691_));
 sky130_fd_sc_hd__nand4_2 _2179_ (.A(_0657_),
    .B(_0670_),
    .C(_0675_),
    .D(_0684_),
    .Y(_0692_));
 sky130_fd_sc_hd__nor2_1 _2180_ (.A(_0659_),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__or2_1 _2181_ (.A(_0659_),
    .B(_0692_),
    .X(_0694_));
 sky130_fd_sc_hd__a22o_1 _2182_ (.A1(\product[46] ),
    .A2(\multiplicand[46] ),
    .B1(\multiplicand[47] ),
    .B2(\product[47] ),
    .X(_0695_));
 sky130_fd_sc_hd__o221a_1 _2183_ (.A1(\product[45] ),
    .A2(\multiplicand[45] ),
    .B1(\multiplicand[46] ),
    .B2(\product[46] ),
    .C1(_0677_),
    .X(_0696_));
 sky130_fd_sc_hd__o22ai_1 _2184_ (.A1(\product[47] ),
    .A2(\multiplicand[47] ),
    .B1(_0695_),
    .B2(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__o221a_2 _2185_ (.A1(_0692_),
    .A2(_0662_),
    .B1(_0627_),
    .B2(_0694_),
    .C1(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__nand2_1 _2186_ (.A(_0628_),
    .B(_0693_),
    .Y(_0699_));
 sky130_fd_sc_hd__o21bai_2 _2187_ (.A1(_0566_),
    .A2(_0559_),
    .B1_N(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__o41a_1 _2188_ (.A1(_0629_),
    .A2(_0659_),
    .A3(_0692_),
    .A4(_0567_),
    .B1(_0698_),
    .X(_0701_));
 sky130_fd_sc_hd__o21ai_4 _2189_ (.A1(_0699_),
    .A2(_0567_),
    .B1(_0698_),
    .Y(_0702_));
 sky130_fd_sc_hd__o21ai_1 _2190_ (.A1(_0691_),
    .A2(_0701_),
    .B1(net133),
    .Y(_0703_));
 sky130_fd_sc_hd__a31o_1 _2191_ (.A1(_0691_),
    .A2(_0698_),
    .A3(_0700_),
    .B1(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__o211a_1 _2192_ (.A1(\product[48] ),
    .A2(net133),
    .B1(_0704_),
    .C1(_0859_),
    .X(_0207_));
 sky130_fd_sc_hd__or2_1 _2193_ (.A(\product[49] ),
    .B(\multiplicand[49] ),
    .X(_0705_));
 sky130_fd_sc_hd__xor2_1 _2194_ (.A(\product[49] ),
    .B(\multiplicand[49] ),
    .X(_0706_));
 sky130_fd_sc_hd__o21a_1 _2195_ (.A1(_0688_),
    .A2(_0701_),
    .B1(_0690_),
    .X(_0707_));
 sky130_fd_sc_hd__o211a_1 _2196_ (.A1(_0688_),
    .A2(_0701_),
    .B1(_0706_),
    .C1(_0690_),
    .X(_0708_));
 sky130_fd_sc_hd__o21ai_1 _2197_ (.A1(_0706_),
    .A2(_0707_),
    .B1(net133),
    .Y(_0709_));
 sky130_fd_sc_hd__o221a_1 _2198_ (.A1(\product[49] ),
    .A2(net133),
    .B1(_0708_),
    .B2(_0709_),
    .C1(_0859_),
    .X(_0208_));
 sky130_fd_sc_hd__nand2_2 _2199_ (.A(\product[50] ),
    .B(\multiplicand[50] ),
    .Y(_0710_));
 sky130_fd_sc_hd__or2_1 _2200_ (.A(\product[50] ),
    .B(\multiplicand[50] ),
    .X(_0711_));
 sky130_fd_sc_hd__nand2_1 _2201_ (.A(_0710_),
    .B(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__and3b_1 _2202_ (.A_N(_0688_),
    .B(_0706_),
    .C(_0690_),
    .X(_0713_));
 sky130_fd_sc_hd__or3b_1 _2203_ (.A(_0688_),
    .B(_0689_),
    .C_N(_0706_),
    .X(_0714_));
 sky130_fd_sc_hd__a22o_1 _2204_ (.A1(\product[48] ),
    .A2(\multiplicand[48] ),
    .B1(\multiplicand[49] ),
    .B2(\product[49] ),
    .X(_0715_));
 sky130_fd_sc_hd__o21ai_1 _2205_ (.A1(\product[49] ),
    .A2(\multiplicand[49] ),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__a22oi_4 _2206_ (.A1(_0705_),
    .A2(_0715_),
    .B1(_0702_),
    .B2(_0713_),
    .Y(_0717_));
 sky130_fd_sc_hd__xnor2_1 _2207_ (.A(_0712_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__a21oi_1 _2208_ (.A1(_0718_),
    .A2(net132),
    .B1(net65),
    .Y(_0719_));
 sky130_fd_sc_hd__o21a_1 _2209_ (.A1(\product[50] ),
    .A2(net132),
    .B1(_0719_),
    .X(_0209_));
 sky130_fd_sc_hd__nor2_1 _2210_ (.A(\product[51] ),
    .B(\multiplicand[51] ),
    .Y(_0720_));
 sky130_fd_sc_hd__or2_2 _2211_ (.A(\product[51] ),
    .B(\multiplicand[51] ),
    .X(_0721_));
 sky130_fd_sc_hd__nand2_1 _2212_ (.A(\product[51] ),
    .B(\multiplicand[51] ),
    .Y(_0722_));
 sky130_fd_sc_hd__o21ai_1 _2213_ (.A1(_0712_),
    .A2(_0717_),
    .B1(_0710_),
    .Y(_0723_));
 sky130_fd_sc_hd__a21boi_1 _2214_ (.A1(_0721_),
    .A2(_0722_),
    .B1_N(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__o2111a_1 _2215_ (.A1(_0712_),
    .A2(_0717_),
    .B1(_0721_),
    .C1(_0722_),
    .D1(_0710_),
    .X(_0725_));
 sky130_fd_sc_hd__a21o_1 _2216_ (.A1(_0844_),
    .A2(\multiplier[0] ),
    .B1(\product[51] ),
    .X(_0726_));
 sky130_fd_sc_hd__o311a_1 _2217_ (.A1(_0725_),
    .A2(_0288_),
    .A3(_0724_),
    .B1(_0726_),
    .C1(_0859_),
    .X(_0210_));
 sky130_fd_sc_hd__nand4_4 _2218_ (.A(_0710_),
    .B(_0711_),
    .C(_0721_),
    .D(_0722_),
    .Y(_0727_));
 sky130_fd_sc_hd__a22oi_4 _2219_ (.A1(\product[50] ),
    .A2(\multiplicand[50] ),
    .B1(\multiplicand[51] ),
    .B2(\product[51] ),
    .Y(_0728_));
 sky130_fd_sc_hd__o22ai_4 _2220_ (.A1(_0720_),
    .A2(_0728_),
    .B1(_0727_),
    .B2(_0717_),
    .Y(_0729_));
 sky130_fd_sc_hd__nand2_1 _2221_ (.A(\product[52] ),
    .B(\multiplicand[52] ),
    .Y(_0730_));
 sky130_fd_sc_hd__or2_1 _2222_ (.A(\product[52] ),
    .B(\multiplicand[52] ),
    .X(_0731_));
 sky130_fd_sc_hd__and2_1 _2223_ (.A(_0730_),
    .B(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__nand2_1 _2224_ (.A(_0729_),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__xnor2_1 _2225_ (.A(_0729_),
    .B(_0732_),
    .Y(_0734_));
 sky130_fd_sc_hd__a21oi_1 _2226_ (.A1(_0844_),
    .A2(\multiplier[0] ),
    .B1(\product[52] ),
    .Y(_0735_));
 sky130_fd_sc_hd__a211oi_1 _2227_ (.A1(_0734_),
    .A2(net132),
    .B1(net65),
    .C1(_0735_),
    .Y(_0211_));
 sky130_fd_sc_hd__or2_1 _2228_ (.A(\product[53] ),
    .B(\multiplicand[53] ),
    .X(_0736_));
 sky130_fd_sc_hd__nand2_1 _2229_ (.A(\product[53] ),
    .B(\multiplicand[53] ),
    .Y(_0737_));
 sky130_fd_sc_hd__a22oi_1 _2230_ (.A1(_0730_),
    .A2(_0733_),
    .B1(_0736_),
    .B2(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__a41o_1 _2231_ (.A1(_0730_),
    .A2(_0733_),
    .A3(_0736_),
    .A4(_0737_),
    .B1(_0288_),
    .X(_0739_));
 sky130_fd_sc_hd__o221a_1 _2232_ (.A1(\product[53] ),
    .A2(net132),
    .B1(_0738_),
    .B2(_0739_),
    .C1(_0859_),
    .X(_0212_));
 sky130_fd_sc_hd__and2_1 _2233_ (.A(\product[54] ),
    .B(\multiplicand[54] ),
    .X(_0740_));
 sky130_fd_sc_hd__nand2_2 _2234_ (.A(\product[54] ),
    .B(\multiplicand[54] ),
    .Y(_0741_));
 sky130_fd_sc_hd__or2_1 _2235_ (.A(\product[54] ),
    .B(\multiplicand[54] ),
    .X(_0742_));
 sky130_fd_sc_hd__and2b_1 _2236_ (.A_N(\product[54] ),
    .B(\multiplicand[54] ),
    .X(_0743_));
 sky130_fd_sc_hd__and2b_1 _2237_ (.A_N(\multiplicand[54] ),
    .B(\product[54] ),
    .X(_0744_));
 sky130_fd_sc_hd__nand2_1 _2238_ (.A(_0741_),
    .B(_0742_),
    .Y(_0745_));
 sky130_fd_sc_hd__a22o_1 _2239_ (.A1(\product[52] ),
    .A2(\multiplicand[52] ),
    .B1(\multiplicand[53] ),
    .B2(\product[53] ),
    .X(_0746_));
 sky130_fd_sc_hd__o21ai_2 _2240_ (.A1(\product[53] ),
    .A2(\multiplicand[53] ),
    .B1(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__and3_1 _2241_ (.A(_0732_),
    .B(_0736_),
    .C(_0737_),
    .X(_0748_));
 sky130_fd_sc_hd__nand2_1 _2242_ (.A(_0729_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__a22oi_1 _2243_ (.A1(_0736_),
    .A2(_0746_),
    .B1(_0729_),
    .B2(_0748_),
    .Y(_0750_));
 sky130_fd_sc_hd__a22oi_1 _2244_ (.A1(_0741_),
    .A2(_0742_),
    .B1(_0729_),
    .B2(_0748_),
    .Y(_0751_));
 sky130_fd_sc_hd__a2bb2oi_1 _2245_ (.A1_N(_0743_),
    .A2_N(_0744_),
    .B1(_0747_),
    .B2(_0749_),
    .Y(_0752_));
 sky130_fd_sc_hd__a21o_1 _2246_ (.A1(_0747_),
    .A2(_0751_),
    .B1(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__o21ai_1 _2247_ (.A1(\product[54] ),
    .A2(net133),
    .B1(_0859_),
    .Y(_0754_));
 sky130_fd_sc_hd__a21oi_1 _2248_ (.A1(_0753_),
    .A2(net133),
    .B1(_0754_),
    .Y(_0213_));
 sky130_fd_sc_hd__xor2_2 _2249_ (.A(\product[55] ),
    .B(\multiplicand[55] ),
    .X(_0755_));
 sky130_fd_sc_hd__o21bai_1 _2250_ (.A1(_0740_),
    .A2(_0752_),
    .B1_N(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__o211ai_1 _2251_ (.A1(_0745_),
    .A2(_0750_),
    .B1(_0755_),
    .C1(_0741_),
    .Y(_0757_));
 sky130_fd_sc_hd__o21ai_1 _2252_ (.A1(\product[55] ),
    .A2(net133),
    .B1(_0859_),
    .Y(_0758_));
 sky130_fd_sc_hd__a31oi_1 _2253_ (.A1(_0756_),
    .A2(_0757_),
    .A3(net133),
    .B1(_0758_),
    .Y(_0214_));
 sky130_fd_sc_hd__nand4_2 _2254_ (.A(_0748_),
    .B(_0755_),
    .C(_0741_),
    .D(_0742_),
    .Y(_0759_));
 sky130_fd_sc_hd__o22a_1 _2255_ (.A1(_0720_),
    .A2(_0728_),
    .B1(_0727_),
    .B2(_0716_),
    .X(_0760_));
 sky130_fd_sc_hd__nor2_1 _2256_ (.A(_0760_),
    .B(_0759_),
    .Y(_0761_));
 sky130_fd_sc_hd__o21ai_1 _2257_ (.A1(\product[55] ),
    .A2(\multiplicand[55] ),
    .B1(_0742_),
    .Y(_0762_));
 sky130_fd_sc_hd__a21oi_1 _2258_ (.A1(_0741_),
    .A2(_0747_),
    .B1(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__a211o_4 _2259_ (.A1(\product[55] ),
    .A2(\multiplicand[55] ),
    .B1(_0761_),
    .C1(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__nor3_1 _2260_ (.A(_0714_),
    .B(_0727_),
    .C(_0759_),
    .Y(_0765_));
 sky130_fd_sc_hd__or3_2 _2261_ (.A(_0714_),
    .B(_0727_),
    .C(_0759_),
    .X(_0766_));
 sky130_fd_sc_hd__a21oi_4 _2262_ (.A1(_0700_),
    .A2(_0698_),
    .B1(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__a21oi_4 _2263_ (.A1(_0702_),
    .A2(_0765_),
    .B1(_0764_),
    .Y(_0768_));
 sky130_fd_sc_hd__and2_1 _2264_ (.A(\product[56] ),
    .B(\multiplicand[56] ),
    .X(_0769_));
 sky130_fd_sc_hd__nor2_1 _2265_ (.A(\product[56] ),
    .B(\multiplicand[56] ),
    .Y(_0770_));
 sky130_fd_sc_hd__or2_1 _2266_ (.A(_0769_),
    .B(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__nor2_1 _2267_ (.A(_0771_),
    .B(_0768_),
    .Y(_0772_));
 sky130_fd_sc_hd__o21a_1 _2268_ (.A1(_0769_),
    .A2(_0770_),
    .B1(_0768_),
    .X(_0773_));
 sky130_fd_sc_hd__nor2_1 _2269_ (.A(_0772_),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__a21o_1 _2270_ (.A1(_0844_),
    .A2(\multiplier[0] ),
    .B1(\product[56] ),
    .X(_0775_));
 sky130_fd_sc_hd__o211a_1 _2271_ (.A1(_0288_),
    .A2(_0774_),
    .B1(_0775_),
    .C1(_0859_),
    .X(_0215_));
 sky130_fd_sc_hd__nor2_1 _2272_ (.A(\product[57] ),
    .B(\multiplicand[57] ),
    .Y(_0776_));
 sky130_fd_sc_hd__and2_1 _2273_ (.A(\product[57] ),
    .B(\multiplicand[57] ),
    .X(_0777_));
 sky130_fd_sc_hd__or2_1 _2274_ (.A(_0776_),
    .B(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__a2111oi_1 _2275_ (.A1(\product[56] ),
    .A2(\multiplicand[56] ),
    .B1(_0772_),
    .C1(_0776_),
    .D1(_0777_),
    .Y(_0779_));
 sky130_fd_sc_hd__o21ai_1 _2276_ (.A1(_0769_),
    .A2(_0772_),
    .B1(_0778_),
    .Y(_0780_));
 sky130_fd_sc_hd__nand2_1 _2277_ (.A(_0780_),
    .B(_0287_),
    .Y(_0781_));
 sky130_fd_sc_hd__o221a_1 _2278_ (.A1(\product[57] ),
    .A2(_0287_),
    .B1(_0779_),
    .B2(_0781_),
    .C1(_0859_),
    .X(_0216_));
 sky130_fd_sc_hd__or2_1 _2279_ (.A(\product[58] ),
    .B(\multiplicand[58] ),
    .X(_0782_));
 sky130_fd_sc_hd__and2_1 _2280_ (.A(\product[58] ),
    .B(\multiplicand[58] ),
    .X(_0783_));
 sky130_fd_sc_hd__nand2_1 _2281_ (.A(\product[58] ),
    .B(\multiplicand[58] ),
    .Y(_0784_));
 sky130_fd_sc_hd__and2_1 _2282_ (.A(_0782_),
    .B(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__nand2_1 _2283_ (.A(_0782_),
    .B(_0784_),
    .Y(_0786_));
 sky130_fd_sc_hd__or4_1 _2284_ (.A(_0769_),
    .B(_0770_),
    .C(_0776_),
    .D(_0777_),
    .X(_0787_));
 sky130_fd_sc_hd__a21oi_1 _2285_ (.A1(\product[57] ),
    .A2(\multiplicand[57] ),
    .B1(_0769_),
    .Y(_0788_));
 sky130_fd_sc_hd__o22ai_2 _2286_ (.A1(_0776_),
    .A2(_0788_),
    .B1(_0787_),
    .B2(_0768_),
    .Y(_0789_));
 sky130_fd_sc_hd__nand2_1 _2287_ (.A(_0789_),
    .B(_0785_),
    .Y(_0790_));
 sky130_fd_sc_hd__xor2_1 _2288_ (.A(_0785_),
    .B(_0789_),
    .X(_0791_));
 sky130_fd_sc_hd__a21o_1 _2289_ (.A1(_0844_),
    .A2(\multiplier[0] ),
    .B1(\product[58] ),
    .X(_0792_));
 sky130_fd_sc_hd__o211a_1 _2290_ (.A1(_0288_),
    .A2(_0791_),
    .B1(_0792_),
    .C1(_0859_),
    .X(_0217_));
 sky130_fd_sc_hd__nor2_1 _2291_ (.A(\product[59] ),
    .B(\multiplicand[59] ),
    .Y(_0793_));
 sky130_fd_sc_hd__and2_1 _2292_ (.A(\product[59] ),
    .B(\multiplicand[59] ),
    .X(_0794_));
 sky130_fd_sc_hd__nand2_1 _2293_ (.A(\product[59] ),
    .B(\multiplicand[59] ),
    .Y(_0795_));
 sky130_fd_sc_hd__nor2_1 _2294_ (.A(_0793_),
    .B(_0794_),
    .Y(_0796_));
 sky130_fd_sc_hd__a21oi_1 _2295_ (.A1(_0784_),
    .A2(_0790_),
    .B1(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__a31o_1 _2296_ (.A1(_0784_),
    .A2(_0790_),
    .A3(_0796_),
    .B1(_0288_),
    .X(_0798_));
 sky130_fd_sc_hd__o221a_1 _2297_ (.A1(\product[59] ),
    .A2(_0287_),
    .B1(_0797_),
    .B2(_0798_),
    .C1(_0859_),
    .X(_0218_));
 sky130_fd_sc_hd__nand2_1 _2298_ (.A(\product[60] ),
    .B(\multiplicand[60] ),
    .Y(_0799_));
 sky130_fd_sc_hd__or2_1 _2299_ (.A(\product[60] ),
    .B(\multiplicand[60] ),
    .X(_0800_));
 sky130_fd_sc_hd__and2_1 _2300_ (.A(_0799_),
    .B(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__o21ai_1 _2301_ (.A1(\product[59] ),
    .A2(\multiplicand[59] ),
    .B1(_0783_),
    .Y(_0802_));
 sky130_fd_sc_hd__or3_1 _2302_ (.A(_0793_),
    .B(_0794_),
    .C(_0786_),
    .X(_0803_));
 sky130_fd_sc_hd__o311a_1 _2303_ (.A1(_0776_),
    .A2(_0788_),
    .A3(_0803_),
    .B1(_0802_),
    .C1(_0795_),
    .X(_0804_));
 sky130_fd_sc_hd__or4_2 _2304_ (.A(_0786_),
    .B(_0793_),
    .C(_0794_),
    .D(_0787_),
    .X(_0805_));
 sky130_fd_sc_hd__o21bai_4 _2305_ (.A1(_0764_),
    .A2(_0767_),
    .B1_N(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__a21bo_1 _2306_ (.A1(_0806_),
    .A2(_0804_),
    .B1_N(_0801_),
    .X(_0807_));
 sky130_fd_sc_hd__o2bb2a_1 _2307_ (.A1_N(_0799_),
    .A2_N(_0800_),
    .B1(_0805_),
    .B2(_0768_),
    .X(_0808_));
 sky130_fd_sc_hd__a21boi_1 _2308_ (.A1(_0804_),
    .A2(_0808_),
    .B1_N(_0807_),
    .Y(_0809_));
 sky130_fd_sc_hd__a21o_1 _2309_ (.A1(_0844_),
    .A2(\multiplier[0] ),
    .B1(\product[60] ),
    .X(_0810_));
 sky130_fd_sc_hd__o211a_1 _2310_ (.A1(_0288_),
    .A2(_0809_),
    .B1(_0810_),
    .C1(_0859_),
    .X(_0219_));
 sky130_fd_sc_hd__nor2_1 _2311_ (.A(\product[61] ),
    .B(\multiplicand[61] ),
    .Y(_0811_));
 sky130_fd_sc_hd__and2_1 _2312_ (.A(\product[61] ),
    .B(\multiplicand[61] ),
    .X(_0812_));
 sky130_fd_sc_hd__nor2_1 _2313_ (.A(_0811_),
    .B(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__a21o_1 _2314_ (.A1(_0799_),
    .A2(_0807_),
    .B1(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__a31oi_1 _2315_ (.A1(_0799_),
    .A2(_0807_),
    .A3(_0813_),
    .B1(_0288_),
    .Y(_0815_));
 sky130_fd_sc_hd__o21ai_1 _2316_ (.A1(\product[61] ),
    .A2(_0287_),
    .B1(_0859_),
    .Y(_0816_));
 sky130_fd_sc_hd__a21oi_1 _2317_ (.A1(_0814_),
    .A2(_0815_),
    .B1(_0816_),
    .Y(_0220_));
 sky130_fd_sc_hd__or2_1 _2318_ (.A(\product[62] ),
    .B(\multiplicand[62] ),
    .X(_0817_));
 sky130_fd_sc_hd__nand2_1 _2319_ (.A(\product[62] ),
    .B(\multiplicand[62] ),
    .Y(_0818_));
 sky130_fd_sc_hd__nand2_1 _2320_ (.A(_0817_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__o21bai_1 _2321_ (.A1(_0799_),
    .A2(_0811_),
    .B1_N(_0812_),
    .Y(_0820_));
 sky130_fd_sc_hd__or3b_1 _2322_ (.A(_0811_),
    .B(_0812_),
    .C_N(_0801_),
    .X(_0821_));
 sky130_fd_sc_hd__a21oi_1 _2323_ (.A1(_0806_),
    .A2(_0804_),
    .B1(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__a21o_1 _2324_ (.A1(_0806_),
    .A2(_0804_),
    .B1(_0821_),
    .X(_0823_));
 sky130_fd_sc_hd__nand3b_1 _2325_ (.A_N(_0820_),
    .B(_0823_),
    .C(_0819_),
    .Y(_0824_));
 sky130_fd_sc_hd__o21bai_2 _2326_ (.A1(_0820_),
    .A2(_0822_),
    .B1_N(_0819_),
    .Y(_0825_));
 sky130_fd_sc_hd__a21oi_1 _2327_ (.A1(_0824_),
    .A2(_0825_),
    .B1(_0288_),
    .Y(_0826_));
 sky130_fd_sc_hd__o21ai_1 _2328_ (.A1(\product[62] ),
    .A2(_0287_),
    .B1(_0859_),
    .Y(_0827_));
 sky130_fd_sc_hd__nor2_1 _2329_ (.A(_0827_),
    .B(_0826_),
    .Y(_0221_));
 sky130_fd_sc_hd__nor2_1 _2330_ (.A(\product[63] ),
    .B(\multiplicand[63] ),
    .Y(_0828_));
 sky130_fd_sc_hd__and2_1 _2331_ (.A(\product[63] ),
    .B(\multiplicand[63] ),
    .X(_0829_));
 sky130_fd_sc_hd__nor2_1 _2332_ (.A(_0828_),
    .B(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__o2bb2ai_1 _2333_ (.A1_N(_0818_),
    .A2_N(_0825_),
    .B1(_0828_),
    .B2(_0829_),
    .Y(_0831_));
 sky130_fd_sc_hd__nand3_1 _2334_ (.A(_0818_),
    .B(_0825_),
    .C(_0830_),
    .Y(_0832_));
 sky130_fd_sc_hd__o21ai_1 _2335_ (.A1(\product[63] ),
    .A2(_0287_),
    .B1(_0859_),
    .Y(_0833_));
 sky130_fd_sc_hd__a31oi_1 _2336_ (.A1(_0831_),
    .A2(_0832_),
    .A3(_0287_),
    .B1(_0833_),
    .Y(_0222_));
 sky130_fd_sc_hd__and4bb_1 _2337_ (.A_N(net24),
    .B_N(_0981_),
    .C(net65),
    .D(net25),
    .X(_0834_));
 sky130_fd_sc_hd__a31o_1 _2338_ (.A1(net140),
    .A2(_0859_),
    .A3(\multiplier[31] ),
    .B1(_0834_),
    .X(_0223_));
 sky130_fd_sc_hd__and2_1 _2339_ (.A(_0844_),
    .B(\count[0] ),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_1 _2340_ (.A(_0859_),
    .B(\count[0] ),
    .Y(_0836_));
 sky130_fd_sc_hd__a21oi_1 _2341_ (.A1(_0867_),
    .A2(_0836_),
    .B1(_0835_),
    .Y(_0224_));
 sky130_fd_sc_hd__and3_1 _2342_ (.A(_0844_),
    .B(\count[1] ),
    .C(\count[0] ),
    .X(_0837_));
 sky130_fd_sc_hd__a21oi_1 _2343_ (.A1(\count[1] ),
    .A2(_0835_),
    .B1(net65),
    .Y(_0838_));
 sky130_fd_sc_hd__o21a_1 _2344_ (.A1(\count[1] ),
    .A2(_0835_),
    .B1(_0838_),
    .X(_0225_));
 sky130_fd_sc_hd__and3_1 _2345_ (.A(\count[2] ),
    .B(\count[1] ),
    .C(_0835_),
    .X(_0839_));
 sky130_fd_sc_hd__a21oi_1 _2346_ (.A1(\count[2] ),
    .A2(_0837_),
    .B1(net65),
    .Y(_0840_));
 sky130_fd_sc_hd__o21a_1 _2347_ (.A1(\count[2] ),
    .A2(_0837_),
    .B1(_0840_),
    .X(_0226_));
 sky130_fd_sc_hd__a31o_1 _2348_ (.A1(\count[3] ),
    .A2(\count[2] ),
    .A3(_0837_),
    .B1(net65),
    .X(_0841_));
 sky130_fd_sc_hd__o21ba_1 _2349_ (.A1(\count[3] ),
    .A2(_0839_),
    .B1_N(_0841_),
    .X(_0227_));
 sky130_fd_sc_hd__a21oi_1 _2350_ (.A1(\count[3] ),
    .A2(_0839_),
    .B1(\count[4] ),
    .Y(_0842_));
 sky130_fd_sc_hd__a311oi_1 _2351_ (.A1(\count[4] ),
    .A2(\count[3] ),
    .A3(_0839_),
    .B1(_0842_),
    .C1(net65),
    .Y(_0228_));
 sky130_fd_sc_hd__and4_1 _2352_ (.A(\count[4] ),
    .B(\count[3] ),
    .C(\count[2] ),
    .D(\count[1] ),
    .X(_0843_));
 sky130_fd_sc_hd__a31o_1 _2353_ (.A1(\count[0] ),
    .A2(_0843_),
    .A3(net142),
    .B1(net136),
    .X(_0229_));
 sky130_fd_sc_hd__dfxtp_4 _2354_ (.CLK(clknet_leaf_20_clk),
    .D(_0000_),
    .Q(\multiplier[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2355_ (.CLK(clknet_leaf_20_clk),
    .D(_0001_),
    .Q(\multiplier[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2356_ (.CLK(clknet_leaf_15_clk),
    .D(_0002_),
    .Q(\multiplier[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2357_ (.CLK(clknet_leaf_15_clk),
    .D(_0003_),
    .Q(\multiplier[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2358_ (.CLK(clknet_leaf_16_clk),
    .D(_0004_),
    .Q(\multiplier[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2359_ (.CLK(clknet_leaf_17_clk),
    .D(_0005_),
    .Q(\multiplier[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2360_ (.CLK(clknet_leaf_16_clk),
    .D(_0006_),
    .Q(\multiplier[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2361_ (.CLK(clknet_leaf_16_clk),
    .D(_0007_),
    .Q(\multiplier[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2362_ (.CLK(clknet_leaf_15_clk),
    .D(_0008_),
    .Q(\multiplier[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2363_ (.CLK(clknet_leaf_15_clk),
    .D(_0009_),
    .Q(\multiplier[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2364_ (.CLK(clknet_leaf_14_clk),
    .D(_0010_),
    .Q(\multiplier[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2365_ (.CLK(clknet_leaf_14_clk),
    .D(_0011_),
    .Q(\multiplier[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2366_ (.CLK(clknet_leaf_13_clk),
    .D(_0012_),
    .Q(\multiplier[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2367_ (.CLK(clknet_leaf_14_clk),
    .D(_0013_),
    .Q(\multiplier[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2368_ (.CLK(clknet_leaf_11_clk),
    .D(_0014_),
    .Q(\multiplier[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2369_ (.CLK(clknet_leaf_10_clk),
    .D(_0015_),
    .Q(\multiplier[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2370_ (.CLK(clknet_leaf_11_clk),
    .D(_0016_),
    .Q(\multiplier[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2371_ (.CLK(clknet_leaf_11_clk),
    .D(_0017_),
    .Q(\multiplier[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2372_ (.CLK(clknet_leaf_11_clk),
    .D(_0018_),
    .Q(\multiplier[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2373_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0019_),
    .Q(\multiplier[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2374_ (.CLK(clknet_leaf_7_clk),
    .D(_0020_),
    .Q(\multiplier[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2375_ (.CLK(clknet_leaf_6_clk),
    .D(_0021_),
    .Q(\multiplier[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2376_ (.CLK(clknet_leaf_6_clk),
    .D(_0022_),
    .Q(\multiplier[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2377_ (.CLK(clknet_leaf_6_clk),
    .D(_0023_),
    .Q(\multiplier[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2378_ (.CLK(clknet_leaf_6_clk),
    .D(_0024_),
    .Q(\multiplier[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2379_ (.CLK(clknet_leaf_5_clk),
    .D(_0025_),
    .Q(\multiplier[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2380_ (.CLK(clknet_leaf_5_clk),
    .D(_0026_),
    .Q(\multiplier[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2381_ (.CLK(clknet_leaf_4_clk),
    .D(_0027_),
    .Q(\multiplier[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2382_ (.CLK(clknet_leaf_4_clk),
    .D(_0028_),
    .Q(\multiplier[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2383_ (.CLK(clknet_leaf_8_clk),
    .D(_0029_),
    .Q(\multiplier[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2384_ (.CLK(clknet_leaf_8_clk),
    .D(_0030_),
    .Q(\multiplier[30] ));
 sky130_fd_sc_hd__dfxtp_2 _2385_ (.CLK(clknet_leaf_1_clk),
    .D(_0031_),
    .Q(\multiplicand[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2386_ (.CLK(clknet_leaf_1_clk),
    .D(_0032_),
    .Q(\multiplicand[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2387_ (.CLK(clknet_leaf_104_clk),
    .D(_0033_),
    .Q(\multiplicand[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2388_ (.CLK(clknet_leaf_104_clk),
    .D(_0034_),
    .Q(\multiplicand[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2389_ (.CLK(clknet_leaf_102_clk),
    .D(_0035_),
    .Q(\multiplicand[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2390_ (.CLK(clknet_leaf_103_clk),
    .D(_0036_),
    .Q(\multiplicand[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2391_ (.CLK(clknet_leaf_101_clk),
    .D(_0037_),
    .Q(\multiplicand[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2392_ (.CLK(clknet_leaf_99_clk),
    .D(_0038_),
    .Q(\multiplicand[7] ));
 sky130_fd_sc_hd__dfxtp_4 _2393_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0039_),
    .Q(\multiplicand[8] ));
 sky130_fd_sc_hd__dfxtp_4 _2394_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0040_),
    .Q(\multiplicand[9] ));
 sky130_fd_sc_hd__dfxtp_2 _2395_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0041_),
    .Q(\multiplicand[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2396_ (.CLK(clknet_leaf_94_clk),
    .D(_0042_),
    .Q(\multiplicand[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2397_ (.CLK(clknet_leaf_94_clk),
    .D(_0043_),
    .Q(\multiplicand[12] ));
 sky130_fd_sc_hd__dfxtp_2 _2398_ (.CLK(clknet_leaf_95_clk),
    .D(_0044_),
    .Q(\multiplicand[13] ));
 sky130_fd_sc_hd__dfxtp_2 _2399_ (.CLK(clknet_leaf_77_clk),
    .D(_0045_),
    .Q(\multiplicand[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2400_ (.CLK(clknet_leaf_76_clk),
    .D(_0046_),
    .Q(\multiplicand[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2401_ (.CLK(clknet_leaf_76_clk),
    .D(_0047_),
    .Q(\multiplicand[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2402_ (.CLK(clknet_leaf_76_clk),
    .D(_0048_),
    .Q(\multiplicand[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2403_ (.CLK(clknet_leaf_75_clk),
    .D(_0049_),
    .Q(\multiplicand[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2404_ (.CLK(clknet_leaf_75_clk),
    .D(_0050_),
    .Q(\multiplicand[19] ));
 sky130_fd_sc_hd__dfxtp_2 _2405_ (.CLK(clknet_leaf_73_clk),
    .D(_0051_),
    .Q(\multiplicand[20] ));
 sky130_fd_sc_hd__dfxtp_2 _2406_ (.CLK(clknet_leaf_70_clk),
    .D(_0052_),
    .Q(\multiplicand[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2407_ (.CLK(clknet_leaf_70_clk),
    .D(_0053_),
    .Q(\multiplicand[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2408_ (.CLK(clknet_leaf_69_clk),
    .D(_0054_),
    .Q(\multiplicand[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2409_ (.CLK(clknet_leaf_69_clk),
    .D(_0055_),
    .Q(\multiplicand[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2410_ (.CLK(clknet_leaf_69_clk),
    .D(_0056_),
    .Q(\multiplicand[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2411_ (.CLK(clknet_leaf_66_clk),
    .D(_0057_),
    .Q(\multiplicand[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2412_ (.CLK(clknet_leaf_83_clk),
    .D(_0058_),
    .Q(\multiplicand[27] ));
 sky130_fd_sc_hd__dfxtp_2 _2413_ (.CLK(clknet_leaf_83_clk),
    .D(_0059_),
    .Q(\multiplicand[28] ));
 sky130_fd_sc_hd__dfxtp_2 _2414_ (.CLK(clknet_leaf_79_clk),
    .D(_0060_),
    .Q(\multiplicand[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2415_ (.CLK(clknet_leaf_79_clk),
    .D(_0061_),
    .Q(\multiplicand[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2416_ (.CLK(clknet_leaf_85_clk),
    .D(_0062_),
    .Q(\multiplicand[31] ));
 sky130_fd_sc_hd__dfxtp_4 _2417_ (.CLK(clknet_leaf_85_clk),
    .D(_0063_),
    .Q(\multiplicand[32] ));
 sky130_fd_sc_hd__dfxtp_1 _2418_ (.CLK(clknet_leaf_62_clk),
    .D(_0064_),
    .Q(\multiplicand[33] ));
 sky130_fd_sc_hd__dfxtp_1 _2419_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0065_),
    .Q(\multiplicand[34] ));
 sky130_fd_sc_hd__dfxtp_1 _2420_ (.CLK(clknet_leaf_61_clk),
    .D(_0066_),
    .Q(\multiplicand[35] ));
 sky130_fd_sc_hd__dfxtp_1 _2421_ (.CLK(clknet_leaf_61_clk),
    .D(_0067_),
    .Q(\multiplicand[36] ));
 sky130_fd_sc_hd__dfxtp_2 _2422_ (.CLK(clknet_leaf_35_clk),
    .D(_0068_),
    .Q(\multiplicand[37] ));
 sky130_fd_sc_hd__dfxtp_1 _2423_ (.CLK(clknet_leaf_36_clk),
    .D(_0069_),
    .Q(\multiplicand[38] ));
 sky130_fd_sc_hd__dfxtp_2 _2424_ (.CLK(clknet_leaf_36_clk),
    .D(_0070_),
    .Q(\multiplicand[39] ));
 sky130_fd_sc_hd__dfxtp_1 _2425_ (.CLK(clknet_leaf_35_clk),
    .D(_0071_),
    .Q(\multiplicand[40] ));
 sky130_fd_sc_hd__dfxtp_2 _2426_ (.CLK(clknet_leaf_34_clk),
    .D(_0072_),
    .Q(\multiplicand[41] ));
 sky130_fd_sc_hd__dfxtp_1 _2427_ (.CLK(clknet_leaf_33_clk),
    .D(_0073_),
    .Q(\multiplicand[42] ));
 sky130_fd_sc_hd__dfxtp_1 _2428_ (.CLK(clknet_leaf_33_clk),
    .D(_0074_),
    .Q(\multiplicand[43] ));
 sky130_fd_sc_hd__dfxtp_2 _2429_ (.CLK(clknet_leaf_33_clk),
    .D(_0075_),
    .Q(\multiplicand[44] ));
 sky130_fd_sc_hd__dfxtp_2 _2430_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0076_),
    .Q(\multiplicand[45] ));
 sky130_fd_sc_hd__dfxtp_2 _2431_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0077_),
    .Q(\multiplicand[46] ));
 sky130_fd_sc_hd__dfxtp_2 _2432_ (.CLK(clknet_leaf_29_clk),
    .D(_0078_),
    .Q(\multiplicand[47] ));
 sky130_fd_sc_hd__dfxtp_1 _2433_ (.CLK(clknet_leaf_37_clk),
    .D(_0079_),
    .Q(\multiplicand[48] ));
 sky130_fd_sc_hd__dfxtp_1 _2434_ (.CLK(clknet_leaf_37_clk),
    .D(_0080_),
    .Q(\multiplicand[49] ));
 sky130_fd_sc_hd__dfxtp_2 _2435_ (.CLK(clknet_leaf_39_clk),
    .D(_0081_),
    .Q(\multiplicand[50] ));
 sky130_fd_sc_hd__dfxtp_2 _2436_ (.CLK(clknet_leaf_39_clk),
    .D(_0082_),
    .Q(\multiplicand[51] ));
 sky130_fd_sc_hd__dfxtp_1 _2437_ (.CLK(clknet_leaf_44_clk),
    .D(_0083_),
    .Q(\multiplicand[52] ));
 sky130_fd_sc_hd__dfxtp_1 _2438_ (.CLK(clknet_leaf_43_clk),
    .D(_0084_),
    .Q(\multiplicand[53] ));
 sky130_fd_sc_hd__dfxtp_2 _2439_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0085_),
    .Q(\multiplicand[54] ));
 sky130_fd_sc_hd__dfxtp_2 _2440_ (.CLK(clknet_leaf_46_clk),
    .D(_0086_),
    .Q(\multiplicand[55] ));
 sky130_fd_sc_hd__dfxtp_4 _2441_ (.CLK(clknet_leaf_47_clk),
    .D(_0087_),
    .Q(\multiplicand[56] ));
 sky130_fd_sc_hd__dfxtp_1 _2442_ (.CLK(clknet_leaf_23_clk),
    .D(_0088_),
    .Q(\multiplicand[57] ));
 sky130_fd_sc_hd__dfxtp_1 _2443_ (.CLK(clknet_leaf_23_clk),
    .D(_0089_),
    .Q(\multiplicand[58] ));
 sky130_fd_sc_hd__dfxtp_1 _2444_ (.CLK(clknet_leaf_24_clk),
    .D(_0090_),
    .Q(\multiplicand[59] ));
 sky130_fd_sc_hd__dfxtp_1 _2445_ (.CLK(clknet_leaf_24_clk),
    .D(_0091_),
    .Q(\multiplicand[60] ));
 sky130_fd_sc_hd__dfxtp_1 _2446_ (.CLK(clknet_leaf_26_clk),
    .D(_0092_),
    .Q(\multiplicand[61] ));
 sky130_fd_sc_hd__dfxtp_1 _2447_ (.CLK(clknet_leaf_26_clk),
    .D(_0093_),
    .Q(\multiplicand[62] ));
 sky130_fd_sc_hd__dfxtp_1 _2448_ (.CLK(clknet_leaf_20_clk),
    .D(_0094_),
    .Q(\multiplicand[63] ));
 sky130_fd_sc_hd__dfxtp_1 _2449_ (.CLK(clknet_leaf_1_clk),
    .D(_0095_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _2450_ (.CLK(clknet_leaf_1_clk),
    .D(_0096_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _2451_ (.CLK(clknet_leaf_0_clk),
    .D(_0097_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _2452_ (.CLK(clknet_leaf_0_clk),
    .D(_0098_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _2453_ (.CLK(clknet_leaf_102_clk),
    .D(_0099_),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_1 _2454_ (.CLK(clknet_leaf_102_clk),
    .D(_0100_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_1 _2455_ (.CLK(clknet_leaf_101_clk),
    .D(_0101_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_1 _2456_ (.CLK(clknet_leaf_100_clk),
    .D(_0102_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_1 _2457_ (.CLK(clknet_leaf_101_clk),
    .D(_0103_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_1 _2458_ (.CLK(clknet_leaf_100_clk),
    .D(_0104_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_4 _2459_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0105_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _2460_ (.CLK(clknet_leaf_95_clk),
    .D(_0106_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _2461_ (.CLK(clknet_leaf_77_clk),
    .D(_0107_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _2462_ (.CLK(clknet_leaf_95_clk),
    .D(_0108_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _2463_ (.CLK(clknet_leaf_77_clk),
    .D(_0109_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _2464_ (.CLK(clknet_leaf_76_clk),
    .D(_0110_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _2465_ (.CLK(clknet_leaf_75_clk),
    .D(_0111_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _2466_ (.CLK(clknet_leaf_75_clk),
    .D(_0112_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _2467_ (.CLK(clknet_leaf_72_clk),
    .D(_0113_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _2468_ (.CLK(clknet_leaf_73_clk),
    .D(_0114_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _2469_ (.CLK(clknet_leaf_71_clk),
    .D(_0115_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _2470_ (.CLK(clknet_leaf_71_clk),
    .D(_0116_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _2471_ (.CLK(clknet_leaf_72_clk),
    .D(_0117_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_1 _2472_ (.CLK(clknet_leaf_71_clk),
    .D(_0118_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _2473_ (.CLK(clknet_leaf_72_clk),
    .D(_0119_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _2474_ (.CLK(clknet_leaf_65_clk),
    .D(_0120_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _2475_ (.CLK(clknet_leaf_71_clk),
    .D(_0121_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_1 _2476_ (.CLK(clknet_leaf_65_clk),
    .D(_0122_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _2477_ (.CLK(clknet_leaf_78_clk),
    .D(_0123_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _2478_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0124_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_1 _2479_ (.CLK(clknet_leaf_77_clk),
    .D(_0125_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _2480_ (.CLK(clknet_leaf_79_clk),
    .D(_0126_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_1 _2481_ (.CLK(clknet_leaf_73_clk),
    .D(_0127_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _2482_ (.CLK(clknet_leaf_54_clk),
    .D(_0128_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_4 _2483_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0129_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _2484_ (.CLK(clknet_leaf_54_clk),
    .D(_0130_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _2485_ (.CLK(clknet_leaf_53_clk),
    .D(_0131_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _2486_ (.CLK(clknet_leaf_53_clk),
    .D(_0132_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _2487_ (.CLK(clknet_leaf_53_clk),
    .D(_0133_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_4 _2488_ (.CLK(clknet_leaf_56_clk),
    .D(_0134_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _2489_ (.CLK(clknet_leaf_76_clk),
    .D(_0135_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _2490_ (.CLK(clknet_leaf_95_clk),
    .D(_0136_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _2491_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0137_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_1 _2492_ (.CLK(clknet_leaf_17_clk),
    .D(_0138_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_1 _2493_ (.CLK(clknet_leaf_17_clk),
    .D(_0139_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_1 _2494_ (.CLK(clknet_leaf_17_clk),
    .D(_0140_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_1 _2495_ (.CLK(clknet_leaf_19_clk),
    .D(_0141_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_1 _2496_ (.CLK(clknet_leaf_19_clk),
    .D(_0142_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_4 _2497_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0143_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_1 _2498_ (.CLK(clknet_leaf_18_clk),
    .D(_0144_),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_1 _2499_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0145_),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_4 _2500_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0146_),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_1 _2501_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0147_),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_4 _2502_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0148_),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_4 _2503_ (.CLK(clknet_leaf_47_clk),
    .D(_0149_),
    .Q(net115));
 sky130_fd_sc_hd__dfxtp_1 _2504_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0150_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_1 _2505_ (.CLK(clknet_leaf_18_clk),
    .D(_0151_),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_1 _2506_ (.CLK(clknet_leaf_18_clk),
    .D(_0152_),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_1 _2507_ (.CLK(clknet_leaf_17_clk),
    .D(_0153_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_1 _2508_ (.CLK(clknet_leaf_17_clk),
    .D(_0154_),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_1 _2509_ (.CLK(clknet_leaf_13_clk),
    .D(_0155_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_1 _2510_ (.CLK(clknet_leaf_10_clk),
    .D(_0156_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_1 _2511_ (.CLK(clknet_leaf_10_clk),
    .D(_0157_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_1 _2512_ (.CLK(clknet_leaf_9_clk),
    .D(_0158_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_4 _2513_ (.CLK(clknet_leaf_1_clk),
    .D(_0159_),
    .Q(\product[0] ));
 sky130_fd_sc_hd__dfxtp_4 _2514_ (.CLK(clknet_leaf_2_clk),
    .D(_0160_),
    .Q(\product[1] ));
 sky130_fd_sc_hd__dfxtp_4 _2515_ (.CLK(clknet_leaf_2_clk),
    .D(_0161_),
    .Q(\product[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2516_ (.CLK(clknet_leaf_103_clk),
    .D(_0162_),
    .Q(\product[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2517_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0163_),
    .Q(\product[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2518_ (.CLK(clknet_leaf_103_clk),
    .D(_0164_),
    .Q(\product[5] ));
 sky130_fd_sc_hd__dfxtp_2 _2519_ (.CLK(clknet_leaf_99_clk),
    .D(_0165_),
    .Q(\product[6] ));
 sky130_fd_sc_hd__dfxtp_2 _2520_ (.CLK(clknet_leaf_99_clk),
    .D(_0166_),
    .Q(\product[7] ));
 sky130_fd_sc_hd__dfxtp_4 _2521_ (.CLK(clknet_leaf_90_clk),
    .D(_0167_),
    .Q(\product[8] ));
 sky130_fd_sc_hd__dfxtp_4 _2522_ (.CLK(clknet_leaf_90_clk),
    .D(_0168_),
    .Q(\product[9] ));
 sky130_fd_sc_hd__dfxtp_4 _2523_ (.CLK(clknet_leaf_92_clk),
    .D(_0169_),
    .Q(\product[10] ));
 sky130_fd_sc_hd__dfxtp_2 _2524_ (.CLK(clknet_leaf_92_clk),
    .D(_0170_),
    .Q(\product[11] ));
 sky130_fd_sc_hd__dfxtp_2 _2525_ (.CLK(clknet_leaf_93_clk),
    .D(_0171_),
    .Q(\product[12] ));
 sky130_fd_sc_hd__dfxtp_4 _2526_ (.CLK(clknet_leaf_93_clk),
    .D(_0172_),
    .Q(\product[13] ));
 sky130_fd_sc_hd__dfxtp_4 _2527_ (.CLK(clknet_leaf_94_clk),
    .D(_0173_),
    .Q(\product[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2528_ (.CLK(clknet_leaf_78_clk),
    .D(_0174_),
    .Q(\product[15] ));
 sky130_fd_sc_hd__dfxtp_2 _2529_ (.CLK(clknet_leaf_78_clk),
    .D(_0175_),
    .Q(\product[16] ));
 sky130_fd_sc_hd__dfxtp_2 _2530_ (.CLK(clknet_leaf_79_clk),
    .D(_0176_),
    .Q(\product[17] ));
 sky130_fd_sc_hd__dfxtp_2 _2531_ (.CLK(clknet_leaf_74_clk),
    .D(_0177_),
    .Q(\product[18] ));
 sky130_fd_sc_hd__dfxtp_2 _2532_ (.CLK(clknet_leaf_74_clk),
    .D(_0178_),
    .Q(\product[19] ));
 sky130_fd_sc_hd__dfxtp_4 _2533_ (.CLK(clknet_leaf_83_clk),
    .D(_0179_),
    .Q(\product[20] ));
 sky130_fd_sc_hd__dfxtp_4 _2534_ (.CLK(clknet_leaf_68_clk),
    .D(_0180_),
    .Q(\product[21] ));
 sky130_fd_sc_hd__dfxtp_2 _2535_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0181_),
    .Q(\product[22] ));
 sky130_fd_sc_hd__dfxtp_2 _2536_ (.CLK(clknet_leaf_68_clk),
    .D(_0182_),
    .Q(\product[23] ));
 sky130_fd_sc_hd__dfxtp_4 _2537_ (.CLK(clknet_leaf_66_clk),
    .D(_0183_),
    .Q(\product[24] ));
 sky130_fd_sc_hd__dfxtp_2 _2538_ (.CLK(clknet_leaf_66_clk),
    .D(_0184_),
    .Q(\product[25] ));
 sky130_fd_sc_hd__dfxtp_2 _2539_ (.CLK(clknet_leaf_84_clk),
    .D(_0185_),
    .Q(\product[26] ));
 sky130_fd_sc_hd__dfxtp_2 _2540_ (.CLK(clknet_leaf_84_clk),
    .D(_0186_),
    .Q(\product[27] ));
 sky130_fd_sc_hd__dfxtp_4 _2541_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0187_),
    .Q(\product[28] ));
 sky130_fd_sc_hd__dfxtp_4 _2542_ (.CLK(clknet_leaf_79_clk),
    .D(_0188_),
    .Q(\product[29] ));
 sky130_fd_sc_hd__dfxtp_2 _2543_ (.CLK(clknet_leaf_81_clk),
    .D(_0189_),
    .Q(\product[30] ));
 sky130_fd_sc_hd__dfxtp_2 _2544_ (.CLK(clknet_leaf_81_clk),
    .D(_0190_),
    .Q(\product[31] ));
 sky130_fd_sc_hd__dfxtp_2 _2545_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0191_),
    .Q(\product[32] ));
 sky130_fd_sc_hd__dfxtp_2 _2546_ (.CLK(clknet_leaf_62_clk),
    .D(_0192_),
    .Q(\product[33] ));
 sky130_fd_sc_hd__dfxtp_2 _2547_ (.CLK(clknet_leaf_60_clk),
    .D(_0193_),
    .Q(\product[34] ));
 sky130_fd_sc_hd__dfxtp_2 _2548_ (.CLK(clknet_leaf_60_clk),
    .D(_0194_),
    .Q(\product[35] ));
 sky130_fd_sc_hd__dfxtp_2 _2549_ (.CLK(clknet_leaf_60_clk),
    .D(_0195_),
    .Q(\product[36] ));
 sky130_fd_sc_hd__dfxtp_2 _2550_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0196_),
    .Q(\product[37] ));
 sky130_fd_sc_hd__dfxtp_2 _2551_ (.CLK(clknet_leaf_56_clk),
    .D(_0197_),
    .Q(\product[38] ));
 sky130_fd_sc_hd__dfxtp_2 _2552_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0198_),
    .Q(\product[39] ));
 sky130_fd_sc_hd__dfxtp_4 _2553_ (.CLK(clknet_leaf_35_clk),
    .D(_0199_),
    .Q(\product[40] ));
 sky130_fd_sc_hd__dfxtp_4 _2554_ (.CLK(clknet_leaf_34_clk),
    .D(_0200_),
    .Q(\product[41] ));
 sky130_fd_sc_hd__dfxtp_2 _2555_ (.CLK(clknet_leaf_34_clk),
    .D(_0201_),
    .Q(\product[42] ));
 sky130_fd_sc_hd__dfxtp_4 _2556_ (.CLK(clknet_leaf_31_clk),
    .D(_0202_),
    .Q(\product[43] ));
 sky130_fd_sc_hd__dfxtp_4 _2557_ (.CLK(clknet_leaf_37_clk),
    .D(_0203_),
    .Q(\product[44] ));
 sky130_fd_sc_hd__dfxtp_4 _2558_ (.CLK(clknet_leaf_31_clk),
    .D(_0204_),
    .Q(\product[45] ));
 sky130_fd_sc_hd__dfxtp_4 _2559_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0205_),
    .Q(\product[46] ));
 sky130_fd_sc_hd__dfxtp_4 _2560_ (.CLK(clknet_leaf_29_clk),
    .D(_0206_),
    .Q(\product[47] ));
 sky130_fd_sc_hd__dfxtp_2 _2561_ (.CLK(clknet_leaf_37_clk),
    .D(_0207_),
    .Q(\product[48] ));
 sky130_fd_sc_hd__dfxtp_2 _2562_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0208_),
    .Q(\product[49] ));
 sky130_fd_sc_hd__dfxtp_4 _2563_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0209_),
    .Q(\product[50] ));
 sky130_fd_sc_hd__dfxtp_4 _2564_ (.CLK(clknet_leaf_39_clk),
    .D(_0210_),
    .Q(\product[51] ));
 sky130_fd_sc_hd__dfxtp_2 _2565_ (.CLK(clknet_leaf_44_clk),
    .D(_0211_),
    .Q(\product[52] ));
 sky130_fd_sc_hd__dfxtp_2 _2566_ (.CLK(clknet_leaf_43_clk),
    .D(_0212_),
    .Q(\product[53] ));
 sky130_fd_sc_hd__dfxtp_2 _2567_ (.CLK(clknet_leaf_46_clk),
    .D(_0213_),
    .Q(\product[54] ));
 sky130_fd_sc_hd__dfxtp_4 _2568_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0214_),
    .Q(\product[55] ));
 sky130_fd_sc_hd__dfxtp_2 _2569_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0215_),
    .Q(\product[56] ));
 sky130_fd_sc_hd__dfxtp_2 _2570_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0216_),
    .Q(\product[57] ));
 sky130_fd_sc_hd__dfxtp_2 _2571_ (.CLK(clknet_leaf_21_clk),
    .D(_0217_),
    .Q(\product[58] ));
 sky130_fd_sc_hd__dfxtp_2 _2572_ (.CLK(clknet_leaf_21_clk),
    .D(_0218_),
    .Q(\product[59] ));
 sky130_fd_sc_hd__dfxtp_2 _2573_ (.CLK(clknet_leaf_26_clk),
    .D(_0219_),
    .Q(\product[60] ));
 sky130_fd_sc_hd__dfxtp_2 _2574_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0220_),
    .Q(\product[61] ));
 sky130_fd_sc_hd__dfxtp_1 _2575_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0221_),
    .Q(\product[62] ));
 sky130_fd_sc_hd__dfxtp_1 _2576_ (.CLK(clknet_leaf_9_clk),
    .D(_0222_),
    .Q(\product[63] ));
 sky130_fd_sc_hd__dfxtp_1 _2577_ (.CLK(clknet_leaf_7_clk),
    .D(_0223_),
    .Q(\multiplier[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2578_ (.CLK(clknet_leaf_87_clk),
    .D(_0224_),
    .Q(\count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2579_ (.CLK(clknet_leaf_87_clk),
    .D(_0225_),
    .Q(\count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2580_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0226_),
    .Q(\count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2581_ (.CLK(clknet_leaf_86_clk),
    .D(_0227_),
    .Q(\count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2582_ (.CLK(clknet_leaf_86_clk),
    .D(_0228_),
    .Q(\count[4] ));
 sky130_fd_sc_hd__dfxtp_4 _2583_ (.CLK(clknet_leaf_86_clk),
    .D(_0229_),
    .Q(\count[5] ));
 sky130_fd_sc_hd__buf_2 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_8 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_16 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_8 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_16 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(b[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_8 input34 (.A(b[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(b[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(b[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(b[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(b[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(b[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(b[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(b[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(b[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(b[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(b[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(b[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(b[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(b[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(b[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(b[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(b[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(b[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(b[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(b[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(b[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(b[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(b[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(b[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(b[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(b[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(b[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(b[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(b[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(b[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(b[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_16 input65 (.A(reset),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_16 output66 (.A(net66),
    .X(mult[0]));
 sky130_fd_sc_hd__clkbuf_16 output67 (.A(net67),
    .X(mult[10]));
 sky130_fd_sc_hd__clkbuf_16 output68 (.A(net68),
    .X(mult[11]));
 sky130_fd_sc_hd__clkbuf_16 output69 (.A(net69),
    .X(mult[12]));
 sky130_fd_sc_hd__clkbuf_16 output70 (.A(net70),
    .X(mult[13]));
 sky130_fd_sc_hd__clkbuf_16 output71 (.A(net71),
    .X(mult[14]));
 sky130_fd_sc_hd__clkbuf_16 output72 (.A(net72),
    .X(mult[15]));
 sky130_fd_sc_hd__clkbuf_16 output73 (.A(net73),
    .X(mult[16]));
 sky130_fd_sc_hd__clkbuf_16 output74 (.A(net74),
    .X(mult[17]));
 sky130_fd_sc_hd__clkbuf_16 output75 (.A(net75),
    .X(mult[18]));
 sky130_fd_sc_hd__clkbuf_16 output76 (.A(net76),
    .X(mult[19]));
 sky130_fd_sc_hd__clkbuf_16 output77 (.A(net77),
    .X(mult[1]));
 sky130_fd_sc_hd__clkbuf_16 output78 (.A(net78),
    .X(mult[20]));
 sky130_fd_sc_hd__clkbuf_16 output79 (.A(net79),
    .X(mult[21]));
 sky130_fd_sc_hd__clkbuf_16 output80 (.A(net80),
    .X(mult[22]));
 sky130_fd_sc_hd__clkbuf_16 output81 (.A(net81),
    .X(mult[23]));
 sky130_fd_sc_hd__clkbuf_16 output82 (.A(net82),
    .X(mult[24]));
 sky130_fd_sc_hd__clkbuf_16 output83 (.A(net83),
    .X(mult[25]));
 sky130_fd_sc_hd__clkbuf_16 output84 (.A(net84),
    .X(mult[26]));
 sky130_fd_sc_hd__clkbuf_16 output85 (.A(net85),
    .X(mult[27]));
 sky130_fd_sc_hd__clkbuf_16 output86 (.A(net86),
    .X(mult[28]));
 sky130_fd_sc_hd__clkbuf_16 output87 (.A(net87),
    .X(mult[29]));
 sky130_fd_sc_hd__clkbuf_16 output88 (.A(net88),
    .X(mult[2]));
 sky130_fd_sc_hd__clkbuf_16 output89 (.A(net89),
    .X(mult[30]));
 sky130_fd_sc_hd__clkbuf_16 output90 (.A(net90),
    .X(mult[31]));
 sky130_fd_sc_hd__clkbuf_16 output91 (.A(net91),
    .X(mult[32]));
 sky130_fd_sc_hd__clkbuf_16 output92 (.A(net92),
    .X(mult[33]));
 sky130_fd_sc_hd__clkbuf_16 output93 (.A(net93),
    .X(mult[34]));
 sky130_fd_sc_hd__clkbuf_16 output94 (.A(net94),
    .X(mult[35]));
 sky130_fd_sc_hd__clkbuf_16 output95 (.A(net95),
    .X(mult[36]));
 sky130_fd_sc_hd__clkbuf_16 output96 (.A(net96),
    .X(mult[37]));
 sky130_fd_sc_hd__clkbuf_16 output97 (.A(net97),
    .X(mult[38]));
 sky130_fd_sc_hd__clkbuf_16 output98 (.A(net98),
    .X(mult[39]));
 sky130_fd_sc_hd__clkbuf_16 output99 (.A(net99),
    .X(mult[3]));
 sky130_fd_sc_hd__clkbuf_16 output100 (.A(net100),
    .X(mult[40]));
 sky130_fd_sc_hd__clkbuf_16 output101 (.A(net101),
    .X(mult[41]));
 sky130_fd_sc_hd__clkbuf_16 output102 (.A(net102),
    .X(mult[42]));
 sky130_fd_sc_hd__clkbuf_16 output103 (.A(net103),
    .X(mult[43]));
 sky130_fd_sc_hd__clkbuf_16 output104 (.A(net104),
    .X(mult[44]));
 sky130_fd_sc_hd__clkbuf_16 output105 (.A(net105),
    .X(mult[45]));
 sky130_fd_sc_hd__clkbuf_16 output106 (.A(net106),
    .X(mult[46]));
 sky130_fd_sc_hd__clkbuf_16 output107 (.A(net107),
    .X(mult[47]));
 sky130_fd_sc_hd__clkbuf_16 output108 (.A(net108),
    .X(mult[48]));
 sky130_fd_sc_hd__clkbuf_16 output109 (.A(net109),
    .X(mult[49]));
 sky130_fd_sc_hd__clkbuf_16 output110 (.A(net110),
    .X(mult[4]));
 sky130_fd_sc_hd__clkbuf_16 output111 (.A(net111),
    .X(mult[50]));
 sky130_fd_sc_hd__clkbuf_16 output112 (.A(net112),
    .X(mult[51]));
 sky130_fd_sc_hd__clkbuf_16 output113 (.A(net113),
    .X(mult[52]));
 sky130_fd_sc_hd__clkbuf_16 output114 (.A(net114),
    .X(mult[53]));
 sky130_fd_sc_hd__clkbuf_16 output115 (.A(net115),
    .X(mult[54]));
 sky130_fd_sc_hd__clkbuf_16 output116 (.A(net116),
    .X(mult[55]));
 sky130_fd_sc_hd__clkbuf_16 output117 (.A(net117),
    .X(mult[56]));
 sky130_fd_sc_hd__clkbuf_16 output118 (.A(net118),
    .X(mult[57]));
 sky130_fd_sc_hd__clkbuf_16 output119 (.A(net119),
    .X(mult[58]));
 sky130_fd_sc_hd__clkbuf_16 output120 (.A(net120),
    .X(mult[59]));
 sky130_fd_sc_hd__clkbuf_16 output121 (.A(net121),
    .X(mult[5]));
 sky130_fd_sc_hd__clkbuf_16 output122 (.A(net122),
    .X(mult[60]));
 sky130_fd_sc_hd__clkbuf_16 output123 (.A(net123),
    .X(mult[61]));
 sky130_fd_sc_hd__clkbuf_16 output124 (.A(net124),
    .X(mult[62]));
 sky130_fd_sc_hd__clkbuf_16 output125 (.A(net125),
    .X(mult[63]));
 sky130_fd_sc_hd__clkbuf_16 output126 (.A(net126),
    .X(mult[6]));
 sky130_fd_sc_hd__clkbuf_16 output127 (.A(net127),
    .X(mult[7]));
 sky130_fd_sc_hd__clkbuf_16 output128 (.A(net128),
    .X(mult[8]));
 sky130_fd_sc_hd__clkbuf_16 output129 (.A(net129),
    .X(mult[9]));
 sky130_fd_sc_hd__buf_8 wire130 (.A(_0350_),
    .X(net130));
 sky130_fd_sc_hd__buf_12 load_slew131 (.A(_0288_),
    .X(net131));
 sky130_fd_sc_hd__buf_12 max_cap132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__buf_12 max_cap133 (.A(_0287_),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_8 max_cap134 (.A(_1153_),
    .X(net134));
 sky130_fd_sc_hd__buf_12 wire135 (.A(_0869_),
    .X(net135));
 sky130_fd_sc_hd__buf_12 max_cap136 (.A(_0869_),
    .X(net136));
 sky130_fd_sc_hd__buf_12 max_cap137 (.A(_0866_),
    .X(net137));
 sky130_fd_sc_hd__buf_12 max_cap138 (.A(_0866_),
    .X(net138));
 sky130_fd_sc_hd__buf_12 max_cap139 (.A(\count[5] ),
    .X(net139));
 sky130_fd_sc_hd__buf_12 max_cap140 (.A(\count[5] ),
    .X(net140));
 sky130_fd_sc_hd__buf_12 max_cap141 (.A(\count[5] ),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_16 load_slew142 (.A(_0859_),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_53_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_54_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_60_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_61_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_62_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_65_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_66_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_68_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_69_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_70_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_71_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_72_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_73_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_74_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_75_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_76_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_77_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_78_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_79_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_81_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_83_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_84_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_85_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_86_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_87_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_90_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_92_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_93_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_94_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_95_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_99_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_100_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_101_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_102_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_103_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_104_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_1_0_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_1_0_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_1_1_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_1_1_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__inv_12 clkload0 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload1 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload2 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__inv_12 clkload3 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload4 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload5 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload6 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload7 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload8 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload9 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload10 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload11 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload12 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload13 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload14 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload15 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload16 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload17 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload18 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload19 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload20 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload21 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload22 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload23 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload24 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload25 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload26 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload27 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload28 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkinv_2 clkload29 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinv_2 clkload30 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__bufinv_16 clkload31 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinv_2 clkload32 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__bufinv_16 clkload33 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__bufinv_16 clkload34 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__bufinv_16 clkload35 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload36 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload37 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload38 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkinv_2 clkload39 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkinv_2 clkload40 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkinv_2 clkload41 (.A(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload42 (.A(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload43 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload44 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkinv_2 clkload45 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload46 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkinv_2 clkload47 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload48 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload49 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload50 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkinv_2 clkload51 (.A(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkinv_2 clkload52 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload53 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkinv_2 clkload54 (.A(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkinv_2 clkload55 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkinv_2 clkload56 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload57 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload58 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkinv_2 clkload59 (.A(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload60 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload61 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload62 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkinv_2 clkload63 (.A(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload64 (.A(clknet_leaf_87_clk));
endmodule
